// Verilog HDL NetList 
//   timeStamp 2009 10 20 10 54 5 
//   author "Avanti Corporation."
//   program "A2Hdl" 
//   design library: cell
//   cell name     : cell.CEL (version 1)
module AFCSHCINX4 ( CI1N , CO0 , S , CO1 , CI0N , CS , A , B );
    input CI1N ;
    output CO0 ;
    output S ;
    output CO1 ;
    input CI0N ;
    input CS ;
    input A ;
    input B ;
endmodule 
module AFCSHCINX2 ( CI1N , CO0 , S , CO1 , CI0N , CS , A , B );
    input CI1N ;
    output CO0 ;
    output S ;
    output CO1 ;
    input CI0N ;
    input CS ;
    input A ;
    input B ;
endmodule 
module ADDHXL ( CO , A , B , S );
    output CO ;
    input A ;
    input B ;
    output S ;
endmodule 
module ADDHX4 ( CO , A , B , S );
    output CO ;
    input A ;
    input B ;
    output S ;
endmodule 
module ADDHX2 ( CO , A , B , S );
    output CO ;
    input A ;
    input B ;
    output S ;
endmodule 
module ADDHX1 ( CO , A , B , S );
    output CO ;
    input A ;
    input B ;
    output S ;
endmodule 
module ADDFXL ( CO , CI , B , A , S );
    output CO ;
    input CI ;
    input B ;
    input A ;
    output S ;
endmodule 
module ADDFX4 ( CO , CI , B , A , S );
    output CO ;
    input CI ;
    input B ;
    input A ;
    output S ;
endmodule 
module ADDFX2 ( CO , CI , B , A , S );
    output CO ;
    input CI ;
    input B ;
    input A ;
    output S ;
endmodule 
module ADDFX1 ( CO , CI , B , A , S );
    output CO ;
    input CI ;
    input B ;
    input A ;
    output S ;
endmodule 
module ADDFHXL ( CO , A , CI , B , S );
    output CO ;
    input A ;
    input CI ;
    input B ;
    output S ;
endmodule 
module ADDFHX4 ( CO , A , CI , B , S );
    output CO ;
    input A ;
    input CI ;
    input B ;
    output S ;
endmodule 
module ADDFHX2 ( CO , A , CI , B , S );
    output CO ;
    input A ;
    input CI ;
    input B ;
    output S ;
endmodule 
module ADDFHX1 ( CO , A , CI , B , S );
    output CO ;
    input A ;
    input CI ;
    input B ;
    output S ;
endmodule 
module AOI21X2 ( B0 , Y , A1 , A0 );
    input B0 ;
    output Y ;
    input A1 ;
    input A0 ;
endmodule 
module AOI21X1 ( B0 , Y , A1 , A0 );
    input B0 ;
    output Y ;
    input A1 ;
    input A0 ;
endmodule 
module AOI211XL ( B0 , Y , C0 , A0 , A1 );
    input B0 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI211X4 ( B0 , Y , C0 , A0 , A1 );
    input B0 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI211X2 ( B0 , Y , C0 , A0 , A1 );
    input B0 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI211X1 ( B0 , Y , C0 , A0 , A1 );
    input B0 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module ANTENNA ( A );
endmodule 
module AND4XL ( D , B , C , A , Y );
    input D ;
    input B ;
    input C ;
    input A ;
    output Y ;
endmodule 
module AND4X4 ( D , B , C , A , Y );
    input D ;
    input B ;
    input C ;
    input A ;
    output Y ;
endmodule 
module AND4X2 ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module AND4X1 ( D , B , C , A , Y );
    input D ;
    input B ;
    input C ;
    input A ;
    output Y ;
endmodule 
module AND3XL ( B , C , A , Y );
    input B ;
    input C ;
    input A ;
    output Y ;
endmodule 
module AND3X4 ( B , C , A , Y );
    input B ;
    input C ;
    input A ;
    output Y ;
endmodule 
module AND3X2 ( B , C , A , Y );
    input B ;
    input C ;
    input A ;
    output Y ;
endmodule 
module AND3X1 ( B , C , A , Y );
    input B ;
    input C ;
    input A ;
    output Y ;
endmodule 
module AND2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AND2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AND2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AND2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AHHCONX4 ( A , CI , S , CON );
    input A ;
    input CI ;
    output S ;
    output CON ;
endmodule 
module AHHCONX2 ( A , CI , S , CON );
    input A ;
    input CI ;
    output S ;
    output CON ;
endmodule 
module AHHCINX4 ( CO , A , CIN , S );
    output CO ;
    input A ;
    input CIN ;
    output S ;
endmodule 
module AHHCINX2 ( CO , A , CIN , S );
    output CO ;
    input A ;
    input CIN ;
    output S ;
endmodule 
module AFHCONX4 ( A , CI , B , S , CON );
    input A ;
    input CI ;
    input B ;
    output S ;
    output CON ;
endmodule 
module AFHCONX2 ( A , CI , B , S , CON );
    input A ;
    input CI ;
    input B ;
    output S ;
    output CON ;
endmodule 
module AFHCINX4 ( CO , A , CIN , B , S );
    output CO ;
    input A ;
    input CIN ;
    input B ;
    output S ;
endmodule 
module AFHCINX2 ( CO , A , CIN , B , S );
    output CO ;
    input A ;
    input CIN ;
    input B ;
    output S ;
endmodule 
module AFCSHCONX4 ( A , B , CO0N , CO1N , S , CS , CI0 , CI1 );
    input A ;
    input B ;
    output CO0N ;
    output CO1N ;
    output S ;
    input CS ;
    input CI0 ;
    input CI1 ;
endmodule 
module AFCSHCONX2 ( A , B , CO0N , CO1N , S , CS , CI0 , CI1 );
    input A ;
    input B ;
    output CO0N ;
    output CO1N ;
    output S ;
    input CS ;
    input CI0 ;
    input CI1 ;
endmodule 
module AOI32X4 ( B0 , B1 , Y , A2 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input A2 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI32X2 ( B1 , B0 , Y , A2 , A0 , A1 );
    input B1 ;
    input B0 ;
    output Y ;
    input A2 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI32X1 ( B0 , B1 , Y , A2 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input A2 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI31XL ( B0 , Y , A2 , A0 , A1 );
    input B0 ;
    output Y ;
    input A2 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI31X4 ( B0 , Y , A2 , A0 , A1 );
    input B0 ;
    output Y ;
    input A2 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI31X2 ( B0 , Y , A0 , A2 , A1 );
    input B0 ;
    output Y ;
    input A0 ;
    input A2 ;
    input A1 ;
endmodule 
module AOI31X1 ( B0 , Y , A2 , A0 , A1 );
    input B0 ;
    output Y ;
    input A2 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI2BB2XL ( B0 , B1 , A0N , Y , A1N );
    input B0 ;
    input B1 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module AOI2BB2X4 ( B0 , B1 , A0N , Y , A1N );
    input B0 ;
    input B1 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module AOI2BB2X2 ( B0 , B1 , A0N , Y , A1N );
    input B0 ;
    input B1 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module AOI2BB2X1 ( B0 , B1 , A0N , Y , A1N );
    input B0 ;
    input B1 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module AOI2BB1XL ( B0 , A0N , Y , A1N );
    input B0 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module AOI2BB1X4 ( B0 , A0N , Y , A1N );
    input B0 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module AOI2BB1X2 ( B0 , A0N , Y , A1N );
    input B0 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module AOI2BB1X1 ( B0 , A0N , Y , A1N );
    input B0 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module AOI22XL ( B1 , B0 , Y , A1 , A0 );
    input B1 ;
    input B0 ;
    output Y ;
    input A1 ;
    input A0 ;
endmodule 
module AOI22X4 ( B1 , B0 , Y , A0 , A1 );
    input B1 ;
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
endmodule 
module AOI22X2 ( B1 , B0 , Y , A1 , A0 );
    input B1 ;
    input B0 ;
    output Y ;
    input A1 ;
    input A0 ;
endmodule 
module AOI22X1 ( B1 , B0 , Y , A1 , A0 );
    input B1 ;
    input B0 ;
    output Y ;
    input A1 ;
    input A0 ;
endmodule 
module AOI222XL ( B0 , B1 , Y , C1 , C0 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input C1 ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI222X4 ( B0 , B1 , Y , C0 , C1 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input C1 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI222X2 ( B0 , B1 , Y , C0 , C1 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input C1 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI222X1 ( B0 , B1 , Y , C1 , C0 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input C1 ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI221XL ( B0 , B1 , Y , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module AOI221X4 ( B0 , B1 , Y , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module AOI221X2 ( B0 , B1 , Y , C0 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module AOI221X1 ( B0 , B1 , Y , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module AOI21XL ( B0 , Y , A1 , A0 );
    input B0 ;
    output Y ;
    input A1 ;
    input A0 ;
endmodule 
module AOI21X4 ( B0 , Y , A1 , A0 );
    input B0 ;
    output Y ;
    input A1 ;
    input A0 ;
endmodule 
module CLKINVX12 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFXL ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX8 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX3 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX2 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX20 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX16 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX12 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFXL ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX8 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX3 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX2 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX20 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX16 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX12 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BMXX1 ( A , M1 , X2 , M0 , S , PP );
    input A ;
    input M1 ;
    input X2 ;
    input M0 ;
    input S ;
    output PP ;
endmodule 
module BENCX4 ( A , M1 , X2 , M2 , M0 , S );
    output A ;
    input M1 ;
    output X2 ;
    input M2 ;
    input M0 ;
    output S ;
endmodule 
module BENCX2 ( A , M1 , X2 , M2 , M0 , S );
    output A ;
    input M1 ;
    output X2 ;
    input M2 ;
    input M0 ;
    output S ;
endmodule 
module BENCX1 ( A , M1 , X2 , M2 , M0 , S );
    output A ;
    input M1 ;
    output X2 ;
    input M2 ;
    input M0 ;
    output S ;
endmodule 
module AOI33XL ( B2 , B0 , B1 , Y , A0 , A1 , A2 );
    input B2 ;
    input B0 ;
    input B1 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module AOI33X4 ( B2 , B0 , B1 , Y , A0 , A1 , A2 );
    input B2 ;
    input B0 ;
    input B1 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module AOI33X2 ( B2 , B0 , B1 , Y , A2 , A1 , A0 );
    input B2 ;
    input B0 ;
    input B1 ;
    output Y ;
    input A2 ;
    input A1 ;
    input A0 ;
endmodule 
module AOI33X1 ( B2 , B0 , B1 , Y , A0 , A1 , A2 );
    input B2 ;
    input B0 ;
    input B1 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module AOI32XL ( B0 , B1 , Y , A2 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input A2 ;
    input A0 ;
    input A1 ;
endmodule 
module DFFNX2 ( CKN , D , QN , Q );
    input CKN ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module DFFNX1 ( CKN , D , QN , Q );
    input CKN ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module DFFNSXL ( CKN , D , SN , QN , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module DFFNSX4 ( CKN , D , SN , QN , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module DFFNSX2 ( CKN , D , SN , QN , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module DFFNSX1 ( CKN , D , SN , QN , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module DFFNSRXL ( CKN , D , SN , QN , RN , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module DFFNSRX4 ( CKN , D , SN , QN , RN , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module DFFNSRX2 ( CKN , D , SN , QN , RN , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module DFFNSRX1 ( CKN , D , SN , QN , RN , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module DFFNRXL ( CKN , D , QN , Q , RN );
    input CKN ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFNRX4 ( CKN , D , QN , Q , RN );
    input CKN ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFNRX2 ( CKN , D , QN , Q , RN );
    input CKN ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFNRX1 ( CKN , D , QN , Q , RN );
    input CKN ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFHQXL ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFHQX4 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFHQX2 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFHQX1 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module CMPR42X2 ( CO , C , B , A , ICO , S , ICI , D );
    output CO ;
    input C ;
    input B ;
    input A ;
    output ICO ;
    output S ;
    input ICI ;
    input D ;
endmodule 
module CMPR42X1 ( CO , C , B , A , ICO , S , ICI , D );
    output CO ;
    input C ;
    input B ;
    input A ;
    output ICO ;
    output S ;
    input ICI ;
    input D ;
endmodule 
module CMPR32X1 ( CO , C , B , A , S );
    output CO ;
    input C ;
    input B ;
    input A ;
    output S ;
endmodule 
module CMPR22X1 ( CO , A , B , S );
    output CO ;
    input A ;
    input B ;
    output S ;
endmodule 
module CLKINVXL ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX8 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX3 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX2 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX20 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX16 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DFFTRX4 ( CK , D , QN , Q , RN );
    input CK ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFTRX2 ( CK , D , QN , Q , RN );
    input CK ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFTRX1 ( CK , D , QN , Q , RN );
    input CK ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFSXL ( CK , D , SN , QN , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module DFFSX4 ( CK , D , SN , QN , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module DFFSX2 ( CK , D , SN , QN , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module DFFSX1 ( CK , D , SN , QN , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module DFFSRXL ( CK , D , SN , QN , RN , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module DFFSRX4 ( CK , D , SN , QN , RN , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module DFFSRX2 ( CK , D , SN , QN , RN , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module DFFSRX1 ( CK , D , SN , QN , RN , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module DFFSRHQXL ( CK , D , SN , RN , Q );
    input CK ;
    input D ;
    input SN ;
    input RN ;
    output Q ;
endmodule 
module DFFSRHQX4 ( CK , D , SN , RN , Q );
    input CK ;
    input D ;
    input SN ;
    input RN ;
    output Q ;
endmodule 
module DFFSRHQX2 ( CK , D , SN , RN , Q );
    input CK ;
    input D ;
    input SN ;
    input RN ;
    output Q ;
endmodule 
module DFFSRHQX1 ( CK , D , SN , RN , Q );
    input CK ;
    input D ;
    input SN ;
    input RN ;
    output Q ;
endmodule 
module DFFSHQXL ( CK , D , SN , Q );
    input CK ;
    input D ;
    input SN ;
    output Q ;
endmodule 
module DFFSHQX4 ( CK , D , SN , Q );
    input CK ;
    input D ;
    input SN ;
    output Q ;
endmodule 
module DFFSHQX2 ( CK , D , SN , Q );
    input CK ;
    input D ;
    input SN ;
    output Q ;
endmodule 
module DFFSHQX1 ( CK , D , SN , Q );
    input CK ;
    input D ;
    input SN ;
    output Q ;
endmodule 
module DFFRXL ( CK , D , QN , Q , RN );
    input CK ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFRX4 ( CK , D , QN , Q , RN );
    input CK ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFRX2 ( CK , D , QN , Q , RN );
    input CK ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFRX1 ( CK , D , QN , Q , RN );
    input CK ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DFFRHQXL ( CK , D , RN , Q );
    input CK ;
    input D ;
    input RN ;
    output Q ;
endmodule 
module DFFRHQX4 ( CK , D , RN , Q );
    input CK ;
    input D ;
    input RN ;
    output Q ;
endmodule 
module DFFRHQX2 ( CK , D , RN , Q );
    input CK ;
    input D ;
    input RN ;
    output Q ;
endmodule 
module DFFRHQX1 ( CK , D , RN , Q );
    input CK ;
    input D ;
    input RN ;
    output Q ;
endmodule 
module DFFNXL ( CKN , D , QN , Q );
    input CKN ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module DFFNX4 ( CKN , D , QN , Q );
    input CKN ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module INVX20 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX16 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX12 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module HOLDX1 ( Y );
    inout Y ;
endmodule 
module FILL8 ();
endmodule 
module FILL64 ();
endmodule 
module FILL4 ();
endmodule 
module FILL32 ();
endmodule 
module FILL2 ();
endmodule 
module FILL16 ();
endmodule 
module FILL1 ();
endmodule 
module EDFFXL ( CK , D , E , QN , Q );
    input CK ;
    input D ;
    input E ;
    output QN ;
    output Q ;
endmodule 
module EDFFX4 ( CK , D , E , QN , Q );
    input CK ;
    input D ;
    input E ;
    output QN ;
    output Q ;
endmodule 
module EDFFX2 ( CK , D , E , QN , Q );
    input CK ;
    input D ;
    input E ;
    output QN ;
    output Q ;
endmodule 
module EDFFX1 ( CK , D , E , QN , Q );
    input CK ;
    input D ;
    input E ;
    output QN ;
    output Q ;
endmodule 
module EDFFTRXL ( CK , D , E , QN , Q , RN );
    input CK ;
    input D ;
    input E ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module EDFFTRX4 ( CK , D , E , QN , Q , RN );
    input CK ;
    input D ;
    input E ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module EDFFTRX2 ( CK , D , E , QN , Q , RN );
    input CK ;
    input D ;
    input E ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module EDFFTRX1 ( CK , D , E , QN , Q , RN );
    input CK ;
    input D ;
    input E ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module DLY4X1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY3X1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY2X1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY1X1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DFFXL ( CK , D , QN , Q );
    input CK ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module DFFX4 ( CK , D , QN , Q );
    input CK ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module DFFX2 ( CK , D , QN , Q );
    input CK ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module DFFX1 ( CK , D , QN , Q );
    input CK ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module DFFTRXL ( CK , D , QN , Q , RN );
    input CK ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module MX4XL ( D , S1 , A , B , C , Y , S0 );
    input D ;
    input S1 ;
    input A ;
    input B ;
    input C ;
    output Y ;
    input S0 ;
endmodule 
module MX4X4 ( D , S0 , S1 , C , A , B , Y );
    input D ;
    input S0 ;
    input S1 ;
    input C ;
    input A ;
    input B ;
    output Y ;
endmodule 
module MX4X2 ( D , S0 , S1 , C , A , B , Y );
    input D ;
    input S0 ;
    input S1 ;
    input C ;
    input A ;
    input B ;
    output Y ;
endmodule 
module MX4X1 ( D , S1 , A , B , C , Y , S0 );
    input D ;
    input S1 ;
    input A ;
    input B ;
    input C ;
    output Y ;
    input S0 ;
endmodule 
module MX2XL ( S0 , B , A , Y );
    input S0 ;
    input B ;
    input A ;
    output Y ;
endmodule 
module MX2X4 ( S0 , B , A , Y );
    input S0 ;
    input B ;
    input A ;
    output Y ;
endmodule 
module MX2X2 ( S0 , B , A , Y );
    input S0 ;
    input B ;
    input A ;
    output Y ;
endmodule 
module MX2X1 ( S0 , B , A , Y );
    input S0 ;
    input B ;
    input A ;
    output Y ;
endmodule 
module JKFFXL ( CK , QN , Q , J , K );
    input CK ;
    output QN ;
    output Q ;
    input J ;
    input K ;
endmodule 
module JKFFX4 ( CK , QN , Q , J , K );
    input CK ;
    output QN ;
    output Q ;
    input J ;
    input K ;
endmodule 
module JKFFX2 ( CK , QN , Q , J , K );
    input CK ;
    output QN ;
    output Q ;
    input J ;
    input K ;
endmodule 
module JKFFX1 ( CK , QN , Q , J , K );
    input CK ;
    output QN ;
    output Q ;
    input J ;
    input K ;
endmodule 
module JKFFSXL ( CK , SN , QN , Q , K , J );
    input CK ;
    input SN ;
    output QN ;
    output Q ;
    input K ;
    input J ;
endmodule 
module JKFFSX4 ( CK , SN , QN , Q , K , J );
    input CK ;
    input SN ;
    output QN ;
    output Q ;
    input K ;
    input J ;
endmodule 
module JKFFSX2 ( CK , SN , QN , Q , K , J );
    input CK ;
    input SN ;
    output QN ;
    output Q ;
    input K ;
    input J ;
endmodule 
module JKFFSX1 ( CK , SN , QN , Q , K , J );
    input CK ;
    input SN ;
    output QN ;
    output Q ;
    input K ;
    input J ;
endmodule 
module JKFFSRXL ( CK , SN , QN , Q , RN , J , K );
    input CK ;
    input SN ;
    output QN ;
    output Q ;
    input RN ;
    input J ;
    input K ;
endmodule 
module JKFFSRX4 ( CK , SN , QN , Q , RN , J , K );
    input CK ;
    input SN ;
    output QN ;
    output Q ;
    input RN ;
    input J ;
    input K ;
endmodule 
module JKFFSRX2 ( CK , SN , QN , Q , RN , J , K );
    input CK ;
    input SN ;
    output QN ;
    output Q ;
    input RN ;
    input J ;
    input K ;
endmodule 
module JKFFSRX1 ( CK , SN , QN , Q , RN , J , K );
    input CK ;
    input SN ;
    output QN ;
    output Q ;
    input RN ;
    input J ;
    input K ;
endmodule 
module JKFFRXL ( CK , QN , Q , RN , K , J );
    input CK ;
    output QN ;
    output Q ;
    input RN ;
    input K ;
    input J ;
endmodule 
module JKFFRX4 ( CK , QN , RN , Q , K , J );
    input CK ;
    output QN ;
    input RN ;
    output Q ;
    input K ;
    input J ;
endmodule 
module JKFFRX2 ( CK , QN , RN , Q , K , J );
    input CK ;
    output QN ;
    input RN ;
    output Q ;
    input K ;
    input J ;
endmodule 
module JKFFRX1 ( CK , QN , Q , RN , K , J );
    input CK ;
    output QN ;
    output Q ;
    input RN ;
    input K ;
    input J ;
endmodule 
module INVXL ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX8 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX3 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX2 ( A , Y );
    input A ;
    output Y ;
endmodule 
module NAND4BX1 ( D , B , AN , C , Y );
    input D ;
    input B ;
    input AN ;
    input C ;
    output Y ;
endmodule 
module NAND4BBXL ( D , AN , C , Y , BN );
    input D ;
    input AN ;
    input C ;
    output Y ;
    input BN ;
endmodule 
module NAND4BBX4 ( D , AN , C , Y , BN );
    input D ;
    input AN ;
    input C ;
    output Y ;
    input BN ;
endmodule 
module NAND4BBX2 ( D , AN , C , Y , BN );
    input D ;
    input AN ;
    input C ;
    output Y ;
    input BN ;
endmodule 
module NAND4BBX1 ( D , AN , C , Y , BN );
    input D ;
    input AN ;
    input C ;
    output Y ;
    input BN ;
endmodule 
module NAND3XL ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NAND3X4 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NAND3X2 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NAND3X1 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NAND3BXL ( C , B , AN , Y );
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NAND3BX4 ( C , B , AN , Y );
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NAND3BX2 ( C , B , AN , Y );
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NAND3BX1 ( C , B , AN , Y );
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NAND2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2BXL ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NAND2BX4 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NAND2BX2 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NAND2BX1 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module MXI4XL ( S0 , S1 , C , A , B , Y , D );
    input S0 ;
    input S1 ;
    input C ;
    input A ;
    input B ;
    output Y ;
    input D ;
endmodule 
module MXI4X4 ( S0 , S1 , C , A , B , Y , D );
    input S0 ;
    input S1 ;
    input C ;
    input A ;
    input B ;
    output Y ;
    input D ;
endmodule 
module MXI4X2 ( S0 , S1 , C , A , B , Y , D );
    input S0 ;
    input S1 ;
    input C ;
    input A ;
    input B ;
    output Y ;
    input D ;
endmodule 
module MXI4X1 ( S0 , S1 , C , A , B , Y , D );
    input S0 ;
    input S1 ;
    input C ;
    input A ;
    input B ;
    output Y ;
    input D ;
endmodule 
module MXI2XL ( S0 , B , A , Y );
    input S0 ;
    input B ;
    input A ;
    output Y ;
endmodule 
module MXI2X4 ( S0 , A , B , Y );
    input S0 ;
    input A ;
    input B ;
    output Y ;
endmodule 
module MXI2X2 ( S0 , B , A , Y );
    input S0 ;
    input B ;
    input A ;
    output Y ;
endmodule 
module MXI2X1 ( S0 , B , A , Y );
    input S0 ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR4BX2 ( D , C , B , AN , Y );
    input D ;
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR4BX1 ( D , C , B , AN , Y );
    input D ;
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR4BBXL ( D , C , AN , Y , BN );
    input D ;
    input C ;
    input AN ;
    output Y ;
    input BN ;
endmodule 
module NOR4BBX4 ( D , C , AN , Y , BN );
    input D ;
    input C ;
    input AN ;
    output Y ;
    input BN ;
endmodule 
module NOR4BBX2 ( D , C , AN , Y , BN );
    input D ;
    input C ;
    input AN ;
    output Y ;
    input BN ;
endmodule 
module NOR4BBX1 ( D , C , AN , Y , BN );
    input D ;
    input C ;
    input AN ;
    output Y ;
    input BN ;
endmodule 
module NOR3XL ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR3X4 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR3X2 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR3X1 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR3BXL ( C , B , AN , Y );
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR3BX4 ( C , B , AN , Y );
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR3BX2 ( C , B , AN , Y );
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR3BX1 ( C , B , AN , Y );
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR2XL ( B , A , Y );
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR2X4 ( B , A , Y );
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR2X2 ( B , A , Y );
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR2X1 ( B , A , Y );
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR2BXL ( B , AN , Y );
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR2BX4 ( B , AN , Y );
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR2BX2 ( B , AN , Y );
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR2BX1 ( B , AN , Y );
    input B ;
    input AN ;
    output Y ;
endmodule 
module NAND4XL ( D , B , A , C , Y );
    input D ;
    input B ;
    input A ;
    input C ;
    output Y ;
endmodule 
module NAND4X4 ( D , B , A , C , Y );
    input D ;
    input B ;
    input A ;
    input C ;
    output Y ;
endmodule 
module NAND4X2 ( D , B , A , C , Y );
    input D ;
    input B ;
    input A ;
    input C ;
    output Y ;
endmodule 
module NAND4X1 ( D , B , A , C , Y );
    input D ;
    input B ;
    input A ;
    input C ;
    output Y ;
endmodule 
module NAND4BXL ( D , B , AN , C , Y );
    input D ;
    input B ;
    input AN ;
    input C ;
    output Y ;
endmodule 
module NAND4BX4 ( D , B , AN , C , Y );
    input D ;
    input B ;
    input AN ;
    input C ;
    output Y ;
endmodule 
module NAND4BX2 ( D , B , AN , C , Y );
    input D ;
    input B ;
    input AN ;
    input C ;
    output Y ;
endmodule 
module OAI2BB1X4 ( B0 , A0N , Y , A1N );
    input B0 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module OAI2BB1X2 ( B0 , A0N , Y , A1N );
    input B0 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module OAI2BB1X1 ( B0 , A0N , Y , A1N );
    input B0 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module OAI22XL ( B0 , B1 , Y , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input A0 ;
    input A1 ;
endmodule 
module OAI22X4 ( B0 , B1 , Y , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input A0 ;
    input A1 ;
endmodule 
module OAI22X2 ( B0 , B1 , Y , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input A1 ;
    input A0 ;
endmodule 
module OAI22X1 ( B0 , B1 , Y , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input A0 ;
    input A1 ;
endmodule 
module OAI222XL ( B0 , B1 , Y , C1 , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C1 ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module OAI222X4 ( B0 , B1 , Y , C1 , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C1 ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module OAI222X2 ( B0 , B1 , Y , C1 , C0 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input C1 ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module OAI222X1 ( B0 , B1 , Y , C1 , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C1 ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module OAI221XL ( B0 , B1 , Y , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module OAI221X4 ( B0 , B1 , Y , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module OAI221X2 ( B0 , B1 , Y , C0 , A0 , A1 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module OAI221X1 ( B0 , B1 , Y , C0 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input C0 ;
    input A1 ;
    input A0 ;
endmodule 
module OAI21XL ( B0 , Y , A0 , A1 );
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
endmodule 
module OAI21X4 ( B0 , Y , A0 , A1 );
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
endmodule 
module OAI21X2 ( B0 , Y , A0 , A1 );
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
endmodule 
module OAI21X1 ( B0 , Y , A0 , A1 );
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
endmodule 
module OAI211XL ( B0 , Y , C0 , A0 , A1 );
    input B0 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module OAI211X4 ( B0 , Y , C0 , A0 , A1 );
    input B0 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module OAI211X2 ( B0 , Y , C0 , A0 , A1 );
    input B0 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module OAI211X1 ( B0 , Y , C0 , A0 , A1 );
    input B0 ;
    output Y ;
    input C0 ;
    input A0 ;
    input A1 ;
endmodule 
module NOR4XL ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR4X4 ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR4X2 ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR4X1 ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module NOR4BXL ( D , C , B , AN , Y );
    input D ;
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module NOR4BX4 ( D , C , B , AN , Y );
    input D ;
    input C ;
    input B ;
    input AN ;
    output Y ;
endmodule 
module OR4XL ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module OR4X4 ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module OR4X2 ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module OR4X1 ( D , C , B , A , Y );
    input D ;
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module OR3XL ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module OR3X4 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module OR3X2 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module OR3X1 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module OR2XL ( B , A , Y );
    input B ;
    input A ;
    output Y ;
endmodule 
module OR2X4 ( B , A , Y );
    input B ;
    input A ;
    output Y ;
endmodule 
module OR2X2 ( B , A , Y );
    input B ;
    input A ;
    output Y ;
endmodule 
module OR2X1 ( B , A , Y );
    input B ;
    input A ;
    output Y ;
endmodule 
module OAI33XL ( B2 , B1 , B0 , Y , A0 , A1 , A2 );
    input B2 ;
    input B1 ;
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module OAI33X4 ( B2 , B1 , B0 , Y , A0 , A1 , A2 );
    input B2 ;
    input B1 ;
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module OAI33X2 ( B2 , B1 , B0 , Y , A1 , A0 , A2 );
    input B2 ;
    input B1 ;
    input B0 ;
    output Y ;
    input A1 ;
    input A0 ;
    input A2 ;
endmodule 
module OAI33X1 ( B2 , B1 , B0 , Y , A0 , A1 , A2 );
    input B2 ;
    input B1 ;
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module OAI32XL ( B0 , B1 , Y , A1 , A2 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input A1 ;
    input A2 ;
    input A0 ;
endmodule 
module OAI32X4 ( B0 , B1 , Y , A2 , A1 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input A2 ;
    input A1 ;
    input A0 ;
endmodule 
module OAI32X2 ( B1 , B0 , Y , A1 , A2 , A0 );
    input B1 ;
    input B0 ;
    output Y ;
    input A1 ;
    input A2 ;
    input A0 ;
endmodule 
module OAI32X1 ( B0 , B1 , Y , A1 , A2 , A0 );
    input B0 ;
    input B1 ;
    output Y ;
    input A1 ;
    input A2 ;
    input A0 ;
endmodule 
module OAI31XL ( B0 , Y , A0 , A1 , A2 );
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module OAI31X4 ( B0 , Y , A2 , A1 , A0 );
    input B0 ;
    output Y ;
    input A2 ;
    input A1 ;
    input A0 ;
endmodule 
module OAI31X2 ( B0 , Y , A0 , A1 , A2 );
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module OAI31X1 ( B0 , Y , A0 , A1 , A2 );
    input B0 ;
    output Y ;
    input A0 ;
    input A1 ;
    input A2 ;
endmodule 
module OAI2BB2XL ( B0 , B1 , Y , A0N , A1N );
    input B0 ;
    input B1 ;
    output Y ;
    input A0N ;
    input A1N ;
endmodule 
module OAI2BB2X4 ( B0 , B1 , Y , A0N , A1N );
    input B0 ;
    input B1 ;
    output Y ;
    input A0N ;
    input A1N ;
endmodule 
module OAI2BB2X2 ( B0 , B1 , Y , A0N , A1N );
    input B0 ;
    input B1 ;
    output Y ;
    input A0N ;
    input A1N ;
endmodule 
module OAI2BB2X1 ( B0 , B1 , Y , A0N , A1N );
    input B0 ;
    input B1 ;
    output Y ;
    input A0N ;
    input A1N ;
endmodule 
module OAI2BB1XL ( B0 , A0N , Y , A1N );
    input B0 ;
    input A0N ;
    output Y ;
    input A1N ;
endmodule 
module SDFFNSXL ( CKN , D , SN , QN , SE , SI , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFNSX4 ( CKN , D , SN , QN , SE , SI , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFNSX2 ( CKN , D , SN , QN , SE , SI , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFNSX1 ( CKN , D , SN , QN , SE , SI , Q );
    input CKN ;
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFNSRXL ( D , SN , QN , SE , SI , RN , Q , CKN );
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
    input CKN ;
endmodule 
module SDFFNSRX4 ( D , SN , QN , SE , SI , RN , Q , CKN );
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
    input CKN ;
endmodule 
module SDFFNSRX2 ( D , SN , QN , SE , SI , RN , Q , CKN );
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
    input CKN ;
endmodule 
module SDFFNSRX1 ( D , SN , QN , SE , SI , RN , Q , CKN );
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
    input CKN ;
endmodule 
module SDFFNRXL ( CKN , D , QN , SE , SI , Q , RN );
    input CKN ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFNRX4 ( CKN , D , QN , SE , SI , Q , RN );
    input CKN ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFNRX2 ( CKN , D , QN , SE , SI , Q , RN );
    input CKN ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFNRX1 ( CKN , D , QN , SE , SI , Q , RN );
    input CKN ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFHQXL ( CK , D , SE , SI , Q );
    input CK ;
    input D ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFHQX4 ( CK , D , SE , SI , Q );
    input CK ;
    input D ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFHQX2 ( CK , D , SE , SI , Q );
    input CK ;
    input D ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFHQX1 ( CK , D , SE , SI , Q );
    input CK ;
    input D ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module RSLATXL ( QN , S , R , Q );
    output QN ;
    input S ;
    input R ;
    output Q ;
endmodule 
module RSLATX4 ( QN , R , S , Q );
    output QN ;
    input R ;
    input S ;
    output Q ;
endmodule 
module RSLATX2 ( QN , R , S , Q );
    output QN ;
    input R ;
    input S ;
    output Q ;
endmodule 
module RSLATX1 ( QN , S , R , Q );
    output QN ;
    input S ;
    input R ;
    output Q ;
endmodule 
module RSLATNXL ( SN , QN , Q , RN );
    input SN ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module RSLATNX4 ( SN , QN , Q , RN );
    input SN ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module RSLATNX2 ( SN , QN , Q , RN );
    input SN ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module RSLATNX1 ( SN , QN , Q , RN );
    input SN ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module RFRDX4 ( RB , BRB );
    input RB ;
    output BRB ;
endmodule 
module RFRDX2 ( RB , BRB );
    input RB ;
    output BRB ;
endmodule 
module RFRDX1 ( RB , BRB );
    input RB ;
    output BRB ;
endmodule 
module RF2R1WX2 ( R1B , R2W , WB , R1W , R2B , WW );
    output R1B ;
    input R2W ;
    input WB ;
    input R1W ;
    output R2B ;
    input WW ;
endmodule 
module RF1R1WX2 ( RB , WB , RW , WW , RWN );
    output RB ;
    input WB ;
    input RW ;
    input WW ;
    input RWN ;
endmodule 
module SDFFTRX1 ( CK , D , QN , SE , SI , Q , RN );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFSXL ( CK , D , SN , QN , SE , SI , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFSX4 ( CK , D , SN , QN , SE , SI , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFSX2 ( CK , D , SN , QN , SE , SI , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFSX1 ( CK , D , SN , QN , SE , SI , Q );
    input CK ;
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFSRXL ( D , SN , QN , SE , SI , RN , Q , CK );
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
    input CK ;
endmodule 
module SDFFSRX4 ( D , SN , QN , SE , SI , RN , Q , CK );
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
    input CK ;
endmodule 
module SDFFSRX2 ( D , SN , QN , SE , SI , RN , Q , CK );
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
    input CK ;
endmodule 
module SDFFSRX1 ( D , SN , QN , SE , SI , RN , Q , CK );
    input D ;
    input SN ;
    output QN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
    input CK ;
endmodule 
module SDFFSRHQXL ( CK , D , SN , SE , SI , RN , Q );
    input CK ;
    input D ;
    input SN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
endmodule 
module SDFFSRHQX4 ( CK , D , SN , SE , SI , RN , Q );
    input CK ;
    input D ;
    input SN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
endmodule 
module SDFFSRHQX2 ( CK , D , SN , SE , SI , RN , Q );
    input CK ;
    input D ;
    input SN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
endmodule 
module SDFFSRHQX1 ( CK , D , SN , SE , SI , RN , Q );
    input CK ;
    input D ;
    input SN ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
endmodule 
module SDFFSHQXL ( CK , D , SN , SE , SI , Q );
    input CK ;
    input D ;
    input SN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFSHQX4 ( CK , D , SN , SE , SI , Q );
    input CK ;
    input D ;
    input SN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFSHQX2 ( CK , D , SN , SE , SI , Q );
    input CK ;
    input D ;
    input SN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFSHQX1 ( CK , D , SN , SE , SI , Q );
    input CK ;
    input D ;
    input SN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFRXL ( CK , D , QN , SE , SI , Q , RN );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFRX4 ( CK , D , QN , SE , SI , Q , RN );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFRX2 ( CK , D , QN , SE , SI , Q , RN );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFRX1 ( CK , D , QN , SE , SI , Q , RN );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFRHQXL ( CK , D , SE , SI , RN , Q );
    input CK ;
    input D ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
endmodule 
module SDFFRHQX4 ( CK , D , SE , SI , RN , Q );
    input CK ;
    input D ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
endmodule 
module SDFFRHQX2 ( CK , D , SE , SI , RN , Q );
    input CK ;
    input D ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
endmodule 
module SDFFRHQX1 ( CK , D , SE , SI , RN , Q );
    input CK ;
    input D ;
    input SE ;
    input SI ;
    input RN ;
    output Q ;
endmodule 
module SDFFNXL ( CKN , D , QN , SE , SI , Q );
    input CKN ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFNX4 ( CKN , D , QN , SE , SI , Q );
    input CKN ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFNX2 ( CKN , D , QN , SE , SI , Q );
    input CKN ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFNX1 ( CKN , D , QN , SE , SI , Q );
    input CKN ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module TBUFX1 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIXL ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIX8 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIX4 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIX3 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIX2 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIX20 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIX16 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIX12 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFIX1 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module SEDFFXL ( CK , D , E , QN , SI , SE , Q );
    input CK ;
    input D ;
    input E ;
    output QN ;
    input SI ;
    input SE ;
    output Q ;
endmodule 
module SEDFFX4 ( CK , D , E , QN , SI , SE , Q );
    input CK ;
    input D ;
    input E ;
    output QN ;
    input SI ;
    input SE ;
    output Q ;
endmodule 
module SEDFFX2 ( CK , D , E , QN , SI , SE , Q );
    input CK ;
    input D ;
    input E ;
    output QN ;
    input SI ;
    input SE ;
    output Q ;
endmodule 
module SEDFFX1 ( CK , D , E , QN , SI , SE , Q );
    input CK ;
    input D ;
    input E ;
    output QN ;
    input SI ;
    input SE ;
    output Q ;
endmodule 
module SEDFFTRXL ( D , E , QN , SI , SE , Q , RN , CK );
    input D ;
    input E ;
    output QN ;
    input SI ;
    input SE ;
    output Q ;
    input RN ;
    input CK ;
endmodule 
module SEDFFTRX4 ( D , E , QN , SI , SE , Q , RN , CK );
    input D ;
    input E ;
    output QN ;
    input SI ;
    input SE ;
    output Q ;
    input RN ;
    input CK ;
endmodule 
module SEDFFTRX2 ( D , E , QN , SI , SE , Q , RN , CK );
    input D ;
    input E ;
    output QN ;
    input SI ;
    input SE ;
    output Q ;
    input RN ;
    input CK ;
endmodule 
module SEDFFTRX1 ( D , E , QN , SI , SE , Q , RN , CK );
    input D ;
    input E ;
    output QN ;
    input SI ;
    input SE ;
    output Q ;
    input RN ;
    input CK ;
endmodule 
module SEDFFHQXL ( CK , D , E , SI , SE , Q );
    input CK ;
    input D ;
    input E ;
    input SI ;
    input SE ;
    output Q ;
endmodule 
module SEDFFHQX4 ( CK , D , E , SI , SE , Q );
    input CK ;
    input D ;
    input E ;
    input SI ;
    input SE ;
    output Q ;
endmodule 
module SEDFFHQX2 ( CK , D , E , SI , SE , Q );
    input CK ;
    input D ;
    input E ;
    input SI ;
    input SE ;
    output Q ;
endmodule 
module SEDFFHQX1 ( CK , D , E , SI , SE , Q );
    input CK ;
    input D ;
    input E ;
    input SI ;
    input SE ;
    output Q ;
endmodule 
module SDFFXL ( CK , D , QN , SE , SI , Q );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFX4 ( CK , D , QN , SE , SI , Q );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFX2 ( CK , D , QN , SE , SI , Q );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFX1 ( CK , D , QN , SE , SI , Q );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
endmodule 
module SDFFTRXL ( CK , D , QN , SE , SI , Q , RN );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFTRX4 ( CK , D , QN , SE , SI , Q , RN );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module SDFFTRX2 ( CK , D , QN , SE , SI , Q , RN );
    input CK ;
    input D ;
    output QN ;
    input SE ;
    input SI ;
    output Q ;
    input RN ;
endmodule 
module TLATRX4 ( D , G , QN , Q , RN );
    input D ;
    input G ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module TLATRX2 ( G , D , QN , Q , RN );
    input G ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module TLATRX1 ( G , D , QN , Q , RN );
    input G ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module TLATNXL ( D , QN , Q , GN );
    input D ;
    output QN ;
    output Q ;
    input GN ;
endmodule 
module TLATNX4 ( D , QN , Q , GN );
    input D ;
    output QN ;
    output Q ;
    input GN ;
endmodule 
module TLATNX2 ( D , QN , Q , GN );
    input D ;
    output QN ;
    output Q ;
    input GN ;
endmodule 
module TLATNX1 ( D , QN , Q , GN );
    input D ;
    output QN ;
    output Q ;
    input GN ;
endmodule 
module TLATNSXL ( D , SN , QN , GN , Q );
    input D ;
    input SN ;
    output QN ;
    input GN ;
    output Q ;
endmodule 
module TLATNSX4 ( D , SN , QN , GN , Q );
    input D ;
    input SN ;
    output QN ;
    input GN ;
    output Q ;
endmodule 
module TLATNSX2 ( D , SN , QN , GN , Q );
    input D ;
    input SN ;
    output QN ;
    input GN ;
    output Q ;
endmodule 
module TLATNSX1 ( D , SN , QN , GN , Q );
    input D ;
    input SN ;
    output QN ;
    input GN ;
    output Q ;
endmodule 
module TLATNSRXL ( D , SN , QN , GN , Q , RN );
    input D ;
    input SN ;
    output QN ;
    input GN ;
    output Q ;
    input RN ;
endmodule 
module TLATNSRX4 ( D , SN , QN , GN , RN , Q );
    input D ;
    input SN ;
    output QN ;
    input GN ;
    input RN ;
    output Q ;
endmodule 
module TLATNSRX2 ( D , SN , QN , GN , Q , RN );
    input D ;
    input SN ;
    output QN ;
    input GN ;
    output Q ;
    input RN ;
endmodule 
module TLATNSRX1 ( D , SN , QN , GN , Q , RN );
    input D ;
    input SN ;
    output QN ;
    input GN ;
    output Q ;
    input RN ;
endmodule 
module TLATNRXL ( D , QN , Q , GN , RN );
    input D ;
    output QN ;
    output Q ;
    input GN ;
    input RN ;
endmodule 
module TLATNRX4 ( D , QN , GN , Q , RN );
    input D ;
    output QN ;
    input GN ;
    output Q ;
    input RN ;
endmodule 
module TLATNRX2 ( D , QN , Q , GN , RN );
    input D ;
    output QN ;
    output Q ;
    input GN ;
    input RN ;
endmodule 
module TLATNRX1 ( D , QN , Q , GN , RN );
    input D ;
    output QN ;
    output Q ;
    input GN ;
    input RN ;
endmodule 
module TIELO ( Y );
    output Y ;
endmodule 
module TIEHI ( Y );
    output Y ;
endmodule 
module TBUFXL ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFX8 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFX4 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFX3 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFX2 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFX20 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFX16 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module TBUFX12 ( A , Y , OE );
    input A ;
    output Y ;
    input OE ;
endmodule 
module XOR3X4 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module XOR3X2 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module XOR2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XOR2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XOR2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XOR2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XNOR3X4 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module XNOR3X2 ( C , B , A , Y );
    input C ;
    input B ;
    input A ;
    output Y ;
endmodule 
module XNOR2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XNOR2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XNOR2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XNOR2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module TTLATXL ( G , D , OE , Q );
    input G ;
    input D ;
    input OE ;
    output Q ;
endmodule 
module TTLATX4 ( D , G , OE , Q );
    input D ;
    input G ;
    input OE ;
    output Q ;
endmodule 
module TTLATX2 ( D , G , OE , Q );
    input D ;
    input G ;
    input OE ;
    output Q ;
endmodule 
module TTLATX1 ( G , D , OE , Q );
    input G ;
    input D ;
    input OE ;
    output Q ;
endmodule 
module TLATXL ( G , D , QN , Q );
    input G ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module TLATX4 ( G , D , QN , Q );
    input G ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module TLATX2 ( G , D , QN , Q );
    input G ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module TLATX1 ( G , D , QN , Q );
    input G ;
    input D ;
    output QN ;
    output Q ;
endmodule 
module TLATSXL ( D , G , SN , QN , Q );
    input D ;
    input G ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module TLATSX4 ( D , G , SN , QN , Q );
    input D ;
    input G ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module TLATSX2 ( D , G , SN , QN , Q );
    input D ;
    input G ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module TLATSX1 ( D , G , SN , QN , Q );
    input D ;
    input G ;
    input SN ;
    output QN ;
    output Q ;
endmodule 
module TLATSRXL ( D , G , SN , QN , Q , RN );
    input D ;
    input G ;
    input SN ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module TLATSRX4 ( G , D , SN , QN , RN , Q );
    input G ;
    input D ;
    input SN ;
    output QN ;
    input RN ;
    output Q ;
endmodule 
module TLATSRX2 ( D , G , SN , QN , Q , RN );
    input D ;
    input G ;
    input SN ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module TLATSRX1 ( D , G , SN , QN , Q , RN );
    input D ;
    input G ;
    input SN ;
    output QN ;
    output Q ;
    input RN ;
endmodule 
module TLATRXL ( G , D , QN , Q , RN );
    input G ;
    input D ;
    output QN ;
    output Q ;
    input RN ;
endmodule 

