* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_shield PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_wos PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT rnod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_s2_std PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_s2_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_s2_sym_ct PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_s3_std PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_s3_sym PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_s3_sym_ct PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT xjvar_nr36 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_w40 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ICV_119
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PDIDGZ C PAD
** N=4 EP=2 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PAD60GU
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PAD60NU
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_118 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X0 1 3 PDIDGZ $T=0 264720 0 270 $X=598 $Y=237040
X1 2 4 PDIDGZ $T=0 344440 0 270 $X=598 $Y=316760
.ENDS
***************************************
.SUBCKT ICV_117 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X0 1 3 PDIDGZ $T=0 424160 0 270 $X=598 $Y=396480
X1 2 4 PDIDGZ $T=0 503880 0 270 $X=598 $Y=476200
.ENDS
***************************************
.SUBCKT ICV_116 2 3 4 5 6 7
** N=11 EP=6 IP=11 FDC=0
X0 2 4 PDIDGZ $T=0 583600 0 270 $X=598 $Y=555920
X1 3 5 PDIDGZ $T=0 663320 0 270 $X=598 $Y=635640
.ENDS
***************************************
.SUBCKT ICV_115 2 3 4 5 6 7
** N=12 EP=6 IP=11 FDC=0
X0 2 4 PDIDGZ $T=0 822760 0 270 $X=598 $Y=795080
X1 3 5 PDIDGZ $T=0 982200 0 270 $X=598 $Y=954520
.ENDS
***************************************
.SUBCKT ICV_114 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X0 1 3 PDIDGZ $T=0 1061920 0 270 $X=598 $Y=1034240
X1 2 4 PDIDGZ $T=0 1141640 0 270 $X=598 $Y=1113960
.ENDS
***************************************
.SUBCKT ICV_113 2 3 4 5 6 7
** N=12 EP=6 IP=11 FDC=0
X0 2 4 PDIDGZ $T=0 1301080 0 270 $X=598 $Y=1273400
X1 3 5 PDIDGZ $T=0 1380800 0 270 $X=598 $Y=1353120
.ENDS
***************************************
.SUBCKT ICV_112 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=15 FDC=0
X0 1 4 PDIDGZ $T=0 1460520 0 270 $X=598 $Y=1432840
X1 3 5 PDIDGZ $T=0 1540240 0 270 $X=598 $Y=1512560
X2 2 6 PDIDGZ $T=0 1619960 0 270 $X=598 $Y=1592280
.ENDS
***************************************
.SUBCKT ICV_111 1 2 3 4
** N=8 EP=4 IP=6 FDC=0
X0 1 2 PDIDGZ $T=0 1779400 0 270 $X=598 $Y=1751720
.ENDS
***************************************
.SUBCKT ICV_110 1 2 3 4
** N=9 EP=4 IP=6 FDC=0
X0 1 2 PDIDGZ $T=0 1938840 0 270 $X=598 $Y=1911160
.ENDS
***************************************
.SUBCKT PDO12CDG I PAD
** N=4 EP=2 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_109 2 3 4 5 6 7
** N=11 EP=6 IP=11 FDC=0
X0 2 4 PDIDGZ $T=0 2018560 0 270 $X=598 $Y=1990880
X4 3 5 PDO12CDG $T=0 2098280 0 270 $X=598 $Y=2070600
.ENDS
***************************************
.SUBCKT ICV_108 2 3 4 5 6 7
** N=12 EP=6 IP=11 FDC=0
X3 2 4 PDO12CDG $T=0 2257720 0 270 $X=598 $Y=2230040
X4 3 5 PDO12CDG $T=0 2417160 0 270 $X=598 $Y=2389480
.ENDS
***************************************
.SUBCKT ICV_107 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X2 2 3 PDO12CDG $T=0 2496880 0 270 $X=598 $Y=2469200
X3 1 4 PDO12CDG $T=0 2576600 0 270 $X=598 $Y=2548920
.ENDS
***************************************
.SUBCKT ICV_106 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=15 FDC=0
X3 1 4 PDO12CDG $T=0 2656320 0 270 $X=598 $Y=2628640
X4 3 6 PDO12CDG $T=0 2736040 0 270 $X=598 $Y=2708360
X5 2 5 PDO12CDG $T=0 2815760 0 270 $X=598 $Y=2788080
.ENDS
***************************************
.SUBCKT ICV_105
** N=6 EP=0 IP=1 FDC=0
.ENDS
***************************************
.SUBCKT ICV_104 1 2 3 4
** N=9 EP=4 IP=6 FDC=0
X2 1 2 PDO12CDG $T=0 2975200 0 270 $X=598 $Y=2947520
.ENDS
***************************************
.SUBCKT ICV_103
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_102 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X2 1 4 PDO12CDG $T=234775 0 0 0 $X=237093 $Y=598
X3 2 3 PDO12CDG $T=314550 0 0 0 $X=316868 $Y=598
.ENDS
***************************************
.SUBCKT ICV_101
** N=2492 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_100
** N=3025 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_99
** N=2406 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_98
** N=3130 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_97
** N=2174 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_96
** N=4108 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_95
** N=2627 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_94
** N=2166 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_93
** N=2844 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_92
** N=3006 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_91
** N=2273 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_90
** N=2318 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX20 A Y VDD VSS
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_89 9 10 12 13 14 233 234
** N=3326 EP=7 IP=12 FDC=0
X0 12 13 10 9 BUFX20 $T=325380 2721040 0 0 $X=325378 $Y=2720638
X1 12 14 10 9 BUFX20 $T=325380 2731120 1 0 $X=325378 $Y=2725680
.ENDS
***************************************
.SUBCKT ICV_88
** N=2050 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_87
** N=2452 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_86 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X0 1 3 PDIDGZ $T=264775 3289640 0 180 $X=237095 $Y=3104640
X1 2 4 PDIDGZ $T=344550 3289640 0 180 $X=316870 $Y=3104640
.ENDS
***************************************
.SUBCKT ICV_85 2 3 4 5 6 7 8 9
** N=13 EP=8 IP=16 FDC=0
X4 2 7 PDO12CDG $T=394325 0 0 0 $X=396643 $Y=598
X5 3 5 PDO12CDG $T=474100 0 0 0 $X=476418 $Y=598
X6 4 6 PDO12CDG $T=633650 0 0 0 $X=635968 $Y=598
.ENDS
***************************************
.SUBCKT ICV_84
** N=4458 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_83
** N=4679 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_82
** N=3780 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_81
** N=5097 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_80
** N=3379 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2X1 B VSS A VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2X4 B VDD VSS A Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2BX1 AN VSS B Y VDD
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI21X1 A1 A0 VSS B0 VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI21XL A1 VSS A0 B0 VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2X4 B A Y VSS VDD
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX1 A VSS VDD Y
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI21X2 A0 A1 VDD B0 Y VSS
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2X1 VDD B A Y VSS
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2X2 A B VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2XL A B VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2X2 A B Y VSS VDD
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI21X4 A0 VDD A1 B0 VSS Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2X2 A VDD B VSS Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2X4 B VSS A VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2X2 A B VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2XL B VSS VDD A Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX4 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI21X1 A1 A0 VDD B0 Y VSS
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI21X2 A1 A0 VSS B0 VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2X4 B A Y VSS VDD
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI21X4 A1 VSS A0 B0 VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX8 A VSS Y VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2X2 B A VDD VSS Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX2 A VSS Y VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_79 2 3 45 47 49 50 51 54 55 56 57 58 59 60 61 62 63 64 65 67
+ 68 69 70 71 73 74 75 76 77 78 79 80 82 84 105 106 136 468 469
** N=6894 EP=39 IP=560 FDC=0
X0 47 3 45 2 1775 NAND2X1 $T=578820 1390480 0 180 $X=576840 $Y=1385040
X1 49 3 50 2 1856 NAND2X1 $T=592680 1390480 0 0 $X=592678 $Y=1390078
X2 54 3 51 2 1886 NAND2X1 $T=599280 1420720 1 180 $X=597300 $Y=1420318
X3 1886 3 1968 2 1970 NAND2X1 $T=605220 1420720 1 0 $X=605218 $Y=1415280
X4 1884 3 1969 2 2004 NAND2X1 $T=605880 1340080 0 0 $X=605878 $Y=1339678
X5 57 3 58 2 1996 NAND2X1 $T=610500 1299760 0 0 $X=610498 $Y=1299358
X6 62 3 60 2 2038 NAND2X1 $T=615780 1319920 0 180 $X=613800 $Y=1314480
X7 2033 3 2059 2 1944 NAND2X1 $T=621060 1390480 1 0 $X=621058 $Y=1385040
X8 65 3 67 2 2089 NAND2X1 $T=625680 1340080 0 0 $X=625678 $Y=1339678
X9 59 3 2120 2 2148 NAND2X1 $T=629640 1420720 0 0 $X=629638 $Y=1420318
X10 2039 3 2216 2 2180 NAND2X1 $T=648120 1269520 1 0 $X=648118 $Y=1264080
X11 47 2 3 45 1826 NOR2X4 $T=587400 1390480 0 180 $X=582780 $Y=1385040
X12 1826 2 3 1860 1973 NOR2X4 $T=598620 1380400 0 0 $X=598618 $Y=1379998
X13 61 2 3 64 2033 NOR2X4 $T=619740 1430800 1 0 $X=619738 $Y=1425360
X14 1826 3 1775 1801 2 NAND2BX1 $T=586740 1380400 1 180 $X=584100 $Y=1379998
X15 1860 3 1856 1857 2 NAND2BX1 $T=595320 1360240 1 180 $X=592680 $Y=1359838
X16 2124 3 2089 2088 2 NAND2BX1 $T=627000 1309840 1 180 $X=624360 $Y=1309438
X17 2160 3 2146 84 2 NAND2BX1 $T=645480 1330000 0 0 $X=645478 $Y=1329598
X18 64 3 59 2222 2 NAND2BX1 $T=650760 1420720 0 0 $X=650758 $Y=1420318
X19 1856 1826 3 1775 2 1829 OAI21X1 $T=593340 1380400 1 180 $X=590040 $Y=1379998
X20 2038 1997 3 1996 2 2098 OAI21X1 $T=619740 1289680 1 0 $X=619738 $Y=1284240
X21 2160 74 3 2146 2 2188 OAI21X1 $T=646140 1319920 1 180 $X=642840 $Y=1319518
X22 1860 3 1858 1856 2 1855 OAI21XL $T=595320 1370320 1 180 $X=592680 $Y=1369918
X23 2180 3 74 2163 2 2151 OAI21XL $T=640860 1259440 0 180 $X=638220 $Y=1254000
X24 2152 3 74 2159 2 2184 OAI21XL $T=644820 1269520 1 180 $X=642180 $Y=1269118
X25 1801 1942 55 3 2 XOR2X4 $T=595320 1350160 0 0 $X=595318 $Y=1349758
X26 2088 2293 105 3 2 XOR2X4 $T=647460 1309840 1 0 $X=647458 $Y=1304400
X27 2222 2161 106 3 2 XOR2X4 $T=647460 1410640 0 0 $X=647458 $Y=1410238
X28 2096 2292 136 3 2 XOR2X4 $T=650760 1259440 0 0 $X=650758 $Y=1259038
X29 1857 3 2 1884 INVX1 $T=595980 1340080 0 0 $X=595978 $Y=1339678
X30 1997 3 2 1976 INVX1 $T=610500 1289680 0 180 $X=609180 $Y=1284240
X31 1858 3 2 2005 INVX1 $T=613800 1370320 1 0 $X=613798 $Y=1364880
X32 2006 3 2 2039 INVX1 $T=614460 1269520 1 0 $X=614458 $Y=1264080
X33 1969 3 2 1971 INVX1 $T=614460 1340080 0 0 $X=614458 $Y=1339678
X34 1944 3 2 2008 INVX1 $T=618420 1370320 0 180 $X=617100 $Y=1364880
X35 2038 3 2 2117 INVX1 $T=619740 1269520 1 0 $X=619738 $Y=1264080
X36 2099 3 2 2159 INVX1 $T=628980 1269520 1 180 $X=627660 $Y=1269118
X37 2216 3 2 2152 INVX1 $T=659340 1269520 0 0 $X=659338 $Y=1269118
X38 56 1943 2 1855 1942 3 AOI21X2 $T=603240 1360240 1 180 $X=598620 $Y=1359838
X39 56 2008 2 2005 1969 3 AOI21X2 $T=616440 1360240 1 180 $X=611820 $Y=1359838
X40 2149 56 2 2151 2123 3 AOI21X2 $T=634920 1239280 0 0 $X=634918 $Y=1238878
X41 2182 56 2 2188 2293 3 AOI21X2 $T=645480 1309840 0 0 $X=645478 $Y=1309438
X42 56 2181 2 2184 2292 3 AOI21X2 $T=654720 1269520 1 180 $X=650100 $Y=1269118
X43 2 1860 1944 1943 3 NOR2X1 $T=601260 1370320 0 0 $X=601258 $Y=1369918
X44 2 2152 73 2181 3 NOR2X1 $T=637560 1269520 0 0 $X=637558 $Y=1269118
X45 2 2160 73 2182 3 NOR2X1 $T=640200 1309840 0 0 $X=640198 $Y=1309438
X46 2 2180 73 2149 3 NOR2X1 $T=642180 1249360 1 180 $X=640200 $Y=1248958
X47 2 64 82 2191 3 NOR2X1 $T=650100 1420720 1 180 $X=648120 $Y=1420318
X48 50 49 3 2 1860 NOR2X2 $T=601260 1390480 0 0 $X=601258 $Y=1390078
X49 58 57 3 2 1997 NOR2X2 $T=609840 1289680 0 0 $X=609838 $Y=1289278
X50 60 62 3 2 2006 NOR2X2 $T=616440 1309840 1 0 $X=616438 $Y=1304400
X51 2006 1997 3 2 2118 NOR2X2 $T=619080 1289680 0 0 $X=619078 $Y=1289278
X52 67 65 3 2 2124 NOR2X2 $T=632940 1340080 0 0 $X=632938 $Y=1339678
X53 2160 2124 3 2 2216 NOR2X2 $T=636900 1299760 0 0 $X=636898 $Y=1299358
X54 77 75 3 2 2160 NOR2X2 $T=643500 1360240 1 0 $X=643498 $Y=1354800
X55 51 54 3 2 1968 OR2XL $T=604560 1420720 0 0 $X=604558 $Y=1420318
X56 1971 1857 1974 3 2 NAND2X2 $T=605880 1340080 1 0 $X=605878 $Y=1334640
X57 77 75 2146 3 2 NAND2X2 $T=638880 1360240 0 180 $X=635580 $Y=1354800
X58 2216 2118 80 3 2 NAND2X2 $T=649440 1289680 0 180 $X=646140 $Y=1284240
X59 1973 2 1999 1829 3 1977 AOI21X4 $T=615120 1380400 1 180 $X=608520 $Y=1379998
X60 2035 2 2033 1999 3 1858 AOI21X4 $T=617760 1390480 1 180 $X=611160 $Y=1390078
X61 2118 2 2099 2098 3 79 AOI21X4 $T=630300 1289680 1 0 $X=630298 $Y=1284240
X62 69 2 2059 2035 3 2161 AOI21X4 $T=632940 1390480 0 0 $X=632938 $Y=1390078
X63 1976 2 1996 3 1998 AND2X2 $T=609840 1279600 1 0 $X=609838 $Y=1274160
X64 1974 3 2004 2 63 NAND2X4 $T=611820 1340080 1 0 $X=611818 $Y=1334640
X65 1886 3 2000 2 1999 NAND2X4 $T=611820 1420720 1 0 $X=611818 $Y=1415280
X66 1973 3 2033 2 71 NAND2X4 $T=622380 1380400 1 0 $X=622378 $Y=1374960
X67 61 59 3 2 2000 OR2X2 $T=615120 1420720 1 180 $X=612480 $Y=1420318
X68 68 64 3 2 2120 OR2X2 $T=637560 1430800 0 180 $X=634920 $Y=1425360
X69 2038 3 2 2039 2096 NAND2XL $T=617100 1259440 0 0 $X=617098 $Y=1259038
X70 68 2035 3 2 INVX4 $T=627000 1390480 1 180 $X=624360 $Y=1390078
X71 2039 2099 2 2117 2163 3 AOI21X1 $T=629640 1259440 0 0 $X=629638 $Y=1259038
X72 2191 69 2 2148 2154 3 AOI21X1 $T=640200 1420720 1 180 $X=637560 $Y=1420318
X73 2146 2124 3 2089 2 2099 OAI21X2 $T=634920 1319920 1 180 $X=629640 $Y=1319518
X74 1998 2123 76 3 2 XNOR2X4 $T=630300 1229200 1 0 $X=630298 $Y=1223760
X75 71 3 68 1977 2 70 OAI21X4 $T=639540 1380400 1 180 $X=632280 $Y=1379998
X76 69 3 56 2 CLKBUFX8 $T=633600 1390480 1 0 $X=633598 $Y=1385040
X77 1970 2154 2 3 78 XOR2X2 $T=635580 1410640 0 0 $X=635578 $Y=1410238
X78 82 3 2059 2 INVX2 $T=653400 1390480 0 0 $X=653398 $Y=1390078
.ENDS
***************************************
.SUBCKT INVXL A VDD VSS Y
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI31X1 A2 A1 A0 VDD B0 Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2X2 B A VDD VSS Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2X1 B A VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2BX1 AN VDD B Y VSS
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDFX2 B A CI CO VDD VSS S
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2X1 B A VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221XL B1 B0 VSS A0 VDD A1 C0 Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDHXL B S A VDD VSS CO
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2XL VDD B A Y VSS
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR3X2 A B C VSS VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI21XL A1 A0 VDD B0 VSS Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB1X1 A1N A0N B0 VSS Y VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_78 1 2 30 32 34 35 36 39 40 41 42 44 45 46 47 48 49 50 51 52
+ 54 55 56 58 59 60 61 62 63 64 65 66 67 68 70 71 72 74 75 76
+ 77 83 84 85 86 87 90 91 92 93 94 95 108 109 110 391 392
** N=4186 EP=57 IP=633 FDC=0
X0 1145 2 30 1 1204 NAND2X1 $T=582120 1521520 1 0 $X=582118 $Y=1516080
X1 1202 2 1189 1 1174 NAND2X1 $T=584760 1521520 1 180 $X=582780 $Y=1521118
X2 1192 2 1203 1 1206 NAND2X1 $T=585420 1582000 1 0 $X=585418 $Y=1576560
X3 1204 2 1190 1 1280 NAND2X1 $T=591360 1481200 1 180 $X=589380 $Y=1480798
X4 47 2 45 1 46 NAND2X1 $T=614460 1440880 0 180 $X=612480 $Y=1435440
X5 1351 2 1336 1 1334 NAND2X1 $T=620400 1481200 1 180 $X=618420 $Y=1480798
X6 1336 2 1358 1 1372 NAND2X1 $T=624360 1481200 0 0 $X=624358 $Y=1480798
X7 1370 2 1337 1 1351 NAND2X1 $T=625680 1551760 1 0 $X=625678 $Y=1546320
X8 1429 2 1431 1 1442 NAND2X1 $T=642840 1501360 0 0 $X=642838 $Y=1500958
X9 1408 2 36 1 1384 NAND2X1 $T=646800 1511440 1 0 $X=646798 $Y=1506000
X10 72 2 74 1 1416 NAND2X1 $T=648120 1461040 1 0 $X=648118 $Y=1455600
X11 39 1 2 40 109 NOR2X4 $T=605220 1430800 0 0 $X=605218 $Y=1430398
X12 72 1 2 74 1428 NOR2X4 $T=648120 1450960 1 0 $X=648118 $Y=1445520
X13 1207 2 1206 1211 1 NAND2BX1 $T=590040 1561840 1 0 $X=590038 $Y=1556400
X14 1428 2 1416 60 1 NAND2BX1 $T=642840 1440880 0 180 $X=640200 $Y=1435440
X15 1317 2 1374 1421 1 NAND2BX1 $T=642840 1531600 1 0 $X=642838 $Y=1526160
X16 1204 1174 2 1209 1 32 OAI21X1 $T=590700 1521520 0 180 $X=587400 $Y=1516080
X17 1173 2 34 1204 1 1223 OAI21XL $T=590040 1471120 0 0 $X=590038 $Y=1470718
X18 1193 2 34 1224 1 1277 OAI21XL $T=591360 1501360 1 0 $X=591358 $Y=1495920
X19 1238 2 34 1229 1 1230 OAI21XL $T=597960 1511440 0 180 $X=595320 $Y=1506000
X20 1350 2 34 1314 1 1312 OAI21XL $T=613800 1471120 1 180 $X=611160 $Y=1470718
X21 1372 2 34 1377 1 1407 OAI21XL $T=627000 1481200 0 0 $X=626998 $Y=1480798
X22 1381 2 1429 1382 1 1356 OAI21XL $T=633600 1511440 1 180 $X=630960 $Y=1511038
X23 86 2 1473 83 1 94 OAI21XL $T=656700 1461040 0 0 $X=656698 $Y=1460638
X24 1206 2 1 1191 INVX1 $T=586080 1561840 0 180 $X=584760 $Y=1556400
X25 1207 2 1 1189 INVX1 $T=587400 1551760 1 180 $X=586080 $Y=1551358
X26 1278 2 1 1205 INVX1 $T=595980 1541680 1 180 $X=594660 $Y=1541278
X27 36 2 1 1238 INVX1 $T=598620 1511440 1 180 $X=597300 $Y=1511038
X28 1282 2 1 1202 INVX1 $T=605220 1531600 1 180 $X=603900 $Y=1531198
X29 1313 2 1 1336 INVX1 $T=611820 1491280 0 0 $X=611818 $Y=1490878
X30 1351 2 1 1368 INVX1 $T=622380 1501360 1 0 $X=622378 $Y=1495920
X31 1356 2 1 1314 INVX1 $T=623700 1471120 1 180 $X=622380 $Y=1470718
X32 61 2 1 1473 INVX1 $T=651420 1461040 0 0 $X=651418 $Y=1460638
X33 1 1145 30 1173 2 NOR2X1 $T=569580 1521520 1 0 $X=569578 $Y=1516080
X34 1 1173 1174 36 2 NOR2X1 $T=577500 1511440 0 0 $X=577498 $Y=1511038
X35 1 1192 1203 1207 2 NOR2X1 $T=585420 1571920 0 0 $X=585418 $Y=1571518
X36 1 1370 1337 1313 2 NOR2X1 $T=620400 1551760 0 180 $X=618420 $Y=1546320
X37 1 1417 1316 1282 2 NOR2X1 $T=620400 1561840 0 180 $X=618420 $Y=1556400
X38 1 1376 54 1381 2 NOR2X1 $T=627000 1511440 1 0 $X=626998 $Y=1506000
X39 1 1381 1384 1358 2 NOR2X1 $T=629640 1501360 1 0 $X=629638 $Y=1495920
X40 1 77 1469 1408 2 NOR2X1 $T=652740 1521520 0 180 $X=650760 $Y=1516080
X41 1 110 63 1469 2 NOR2X1 $T=661980 1541680 0 180 $X=660000 $Y=1536240
X42 45 47 2 1 51 NOR2X2 $T=619740 1440880 1 0 $X=619738 $Y=1435440
X43 86 1428 2 1 62 NOR2X2 $T=655380 1450960 0 0 $X=655378 $Y=1450558
X44 87 92 2 1 86 NOR2X2 $T=659340 1481200 0 180 $X=656040 $Y=1475760
X45 1419 1416 1411 2 1 NAND2X2 $T=639540 1440880 0 0 $X=639538 $Y=1440478
X46 87 92 83 2 1 NAND2X2 $T=658020 1481200 0 0 $X=658018 $Y=1480798
X47 62 1 61 1411 2 59 AOI21X4 $T=644160 1450960 1 180 $X=637560 $Y=1450558
X48 1313 1317 2 1 1347 OR2X2 $T=613800 1531600 1 0 $X=613798 $Y=1526160
X49 34 1384 2 1 1431 OR2X2 $T=634920 1501360 0 0 $X=634918 $Y=1500958
X50 1428 83 2 1 1419 OR2X2 $T=654060 1440880 0 0 $X=654058 $Y=1440478
X51 1189 2 1 1190 1193 NAND2XL $T=584100 1501360 1 0 $X=584098 $Y=1495920
X52 1417 2 1 1316 1278 NAND2XL $T=610500 1561840 0 180 $X=608520 $Y=1556400
X53 56 2 1 1391 1374 NAND2XL $T=631620 1541680 0 180 $X=629640 $Y=1536240
X54 1376 2 1 54 1382 NAND2XL $T=634260 1521520 0 180 $X=632280 $Y=1516080
X55 1406 2 1 1408 64 NAND2XL $T=637560 1521520 1 0 $X=637558 $Y=1516080
X56 1191 1202 1 1205 1209 2 AOI21X1 $T=585420 1541680 1 0 $X=585418 $Y=1536240
X57 1356 1336 1 1368 1377 2 AOI21X1 $T=624360 1491280 1 0 $X=624358 $Y=1485840
X58 1408 32 1 66 1429 2 AOI21X1 $T=646800 1521520 0 180 $X=644160 $Y=1516080
X59 1281 1277 1 2 41 XOR2X2 $T=601260 1501360 1 0 $X=601258 $Y=1495920
X60 1173 1 2 1190 INVXL $T=580140 1481200 0 0 $X=580138 $Y=1480798
X61 32 1 2 1229 INVXL $T=592020 1511440 0 180 $X=590700 $Y=1506000
X62 1358 1 2 1350 INVXL $T=631620 1471120 1 180 $X=630300 $Y=1470718
X63 1469 1 2 108 INVXL $T=660000 1511440 0 0 $X=659998 $Y=1511038
X64 1145 30 1189 1 1191 1224 2 AOI31X1 $T=586080 1531600 1 0 $X=586078 $Y=1526160
X65 1211 1223 1 2 35 XNOR2X2 $T=588060 1461040 0 0 $X=588058 $Y=1460638
X66 48 1230 1 2 42 XNOR2X2 $T=616440 1511440 0 180 $X=609180 $Y=1506000
X67 34 1280 2 1 44 XOR2X1 $T=600600 1471120 0 0 $X=600598 $Y=1470718
X68 1278 1 1282 1281 2 NOR2BX1 $T=607200 1541680 1 180 $X=604560 $Y=1541278
X69 1413 52 49 1203 1 2 1145 ADDFX2 $T=628320 1592080 1 180 $X=614460 $Y=1591678
X70 1414 1371 1348 1316 1 2 1192 ADDFX2 $T=630300 1582000 1 180 $X=616440 $Y=1581598
X71 93 55 65 1423 1 2 1371 ADDFX2 $T=652740 1571920 1 180 $X=638880 $Y=1571518
X72 67 58 55 1425 1 2 1418 ADDFX2 $T=653400 1592080 0 180 $X=639540 $Y=1586640
X73 85 1468 1418 1348 1 2 1413 ADDFX2 $T=654060 1592080 1 180 $X=640200 $Y=1591678
X74 84 1423 1430 63 1 2 1417 ADDFX2 $T=654720 1561840 1 180 $X=640860 $Y=1561438
X75 1471 56 1425 1430 1 2 1414 ADDFX2 $T=654720 1582000 0 180 $X=640860 $Y=1576560
X76 1334 1312 2 1 50 XNOR2X1 $T=616440 1461040 1 0 $X=616438 $Y=1455600
X77 1421 1407 2 1 68 XNOR2X1 $T=640200 1481200 0 0 $X=640198 $Y=1480798
X78 1347 1382 2 1317 1 1351 1374 1378 OAI221XL $T=629640 1531600 0 180 $X=625020 $Y=1526160
X79 58 1370 55 1 2 1391 ADDHXL $T=639540 1551760 1 180 $X=632280 $Y=1551358
X80 70 1376 67 1 2 1337 ADDHXL $T=650760 1551760 0 180 $X=643500 $Y=1546320
X81 71 1468 75 1 2 1471 ADDHXL $T=645480 1602160 0 0 $X=645478 $Y=1601758
X82 1 1381 1347 1406 2 NOR2XL $T=634920 1531600 1 0 $X=634918 $Y=1526160
X83 1 56 1391 1317 2 NOR2XL $T=636240 1541680 0 0 $X=636238 $Y=1541278
X84 54 1376 1442 2 1 76 XOR3X2 $T=638220 1491280 0 0 $X=638218 $Y=1490878
X85 1406 66 1 1378 2 91 AOI21XL $T=654720 1521520 0 0 $X=654718 $Y=1521118
X86 108 32 95 2 90 1 OAI2BB1X1 $T=661320 1511440 0 180 $X=658020 $Y=1506000
.ENDS
***************************************
.SUBCKT NAND2BXL AN VSS B VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX3 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB2X1 A1N A0N B1 B0 VDD VSS Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDFHX1 A B CI CO VDD VSS S
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3X1 C VSS B VDD A Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CMPR32X1 B A C CO VSS VDD S
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_77 1 3 16 17 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34
+ 35 36 37 38 39 40 41 42 43 44 45 46 47 48 50 51 52 53 54 61
+ 63 75 344 345
** N=3605 EP=44 IP=604 FDC=0
X0 1067 1 1064 3 1033 NAND2X1 $T=571560 1733200 0 180 $X=569580 $Y=1727760
X1 28 1 1079 3 1049 NAND2X1 $T=576840 1763440 1 180 $X=574860 $Y=1763038
X2 1120 1 1098 3 937 NAND2X1 $T=590700 1702960 1 0 $X=590698 $Y=1697520
X3 1173 1 1122 3 1062 NAND2X1 $T=599940 1662640 0 0 $X=599938 $Y=1662238
X4 1191 1 1190 3 1189 NAND2X1 $T=607860 1723120 0 180 $X=605880 $Y=1717680
X5 1205 1 1190 3 1192 NAND2X1 $T=611160 1723120 0 180 $X=609180 $Y=1717680
X6 1191 1 1205 3 1188 NAND2X1 $T=611820 1713040 1 0 $X=611818 $Y=1707600
X7 1045 1 1049 1019 3 NAND2BX1 $T=569580 1773520 0 180 $X=566940 $Y=1768080
X8 1033 939 1 937 3 1016 OAI21X1 $T=562320 1702960 0 180 $X=559020 $Y=1697520
X9 1007 997 1 1063 3 1066 OAI21X1 $T=572880 1692880 0 180 $X=569580 $Y=1687440
X10 957 1 19 1007 3 1018 OAI21XL $T=554400 1733200 0 0 $X=554398 $Y=1732798
X11 1034 1 1069 1062 3 958 OAI21XL $T=572220 1672720 1 0 $X=572218 $Y=1667280
X12 1062 1 1101 1095 3 1065 OAI21XL $T=586740 1652560 1 180 $X=584100 $Y=1652158
X13 1007 1 3 959 INVX1 $T=547800 1682800 0 180 $X=546480 $Y=1677360
X14 24 1 3 25 INVX1 $T=564300 1773520 0 0 $X=564298 $Y=1773118
X15 1016 1 3 1069 INVX1 $T=567600 1672720 1 0 $X=567598 $Y=1667280
X16 1015 24 3 1044 1007 1 AOI21X2 $T=562320 1753360 0 0 $X=562318 $Y=1752958
X17 3 1045 21 1015 1 NOR2X1 $T=557700 1773520 0 180 $X=555720 $Y=1768080
X18 3 28 1079 1045 1 NOR2X1 $T=576840 1773520 1 180 $X=574860 $Y=1773118
X19 3 1101 1034 1043 1 NOR2X1 $T=578820 1662640 1 180 $X=576840 $Y=1662238
X20 3 1173 1122 1034 1 NOR2X1 $T=593340 1662640 1 180 $X=591360 $Y=1662238
X21 3 1175 1129 1101 1 NOR2X1 $T=596640 1652560 0 180 $X=594660 $Y=1647120
X22 957 997 1 3 960 NOR2X2 $T=549120 1692880 0 180 $X=545820 $Y=1687440
X23 1001 939 1 3 1003 NOR2X2 $T=548460 1702960 1 0 $X=548458 $Y=1697520
X24 1064 1067 1 3 1001 NOR2X2 $T=579480 1723120 1 0 $X=579478 $Y=1717680
X25 1098 1120 1 3 939 NOR2X2 $T=584100 1702960 0 180 $X=580800 $Y=1697520
X26 20 1015 957 1 3 NAND2X2 $T=556380 1753360 1 180 $X=553080 $Y=1752958
X27 1043 1003 997 1 3 NAND2X2 $T=563640 1672720 0 0 $X=563638 $Y=1672318
X28 938 3 960 1066 1 31 AOI21X4 $T=578820 1692880 1 0 $X=578818 $Y=1687440
X29 955 3 936 1 922 AND2X2 $T=535260 1672720 0 180 $X=532620 $Y=1667280
X30 936 3 1003 1 1005 AND2X2 $T=551100 1672720 1 0 $X=551098 $Y=1667280
X31 1079 28 1 3 1093 OR2X2 $T=592680 1773520 0 180 $X=590040 $Y=1768080
X32 1175 1 3 1129 1095 NAND2XL $T=601920 1642480 1 180 $X=599940 $Y=1642078
X33 16 19 1 3 INVX4 $T=548460 1753360 1 180 $X=545820 $Y=1752958
X34 955 959 3 958 941 1 AOI21X1 $T=547140 1672720 0 180 $X=544500 $Y=1667280
X35 1003 959 3 1016 1006 1 AOI21X1 $T=555060 1682800 1 0 $X=555058 $Y=1677360
X36 1016 1043 3 1065 1063 1 AOI21X1 $T=569580 1672720 0 0 $X=569578 $Y=1672318
X37 908 923 17 1 3 XNOR2X4 $T=530640 1692880 0 0 $X=530638 $Y=1692478
X38 1019 22 27 1 3 XNOR2X4 $T=559020 1763440 0 0 $X=559018 $Y=1763038
X39 957 3 1 936 INVXL $T=539880 1692880 0 180 $X=538560 $Y=1687440
X40 1017 1018 3 1 23 XNOR2X2 $T=555720 1723120 0 0 $X=555718 $Y=1722718
X41 1050 1048 3 1 26 XNOR2X2 $T=567600 1632400 1 0 $X=567598 $Y=1626960
X42 1080 956 3 1 29 XNOR2X2 $T=575520 1642480 1 0 $X=575518 $Y=1637040
X43 1190 1205 1 3 1218 XOR2X1 $T=613800 1723120 1 0 $X=613798 $Y=1717680
X44 1218 1191 1 3 1110 XOR2X1 $T=619080 1723120 1 180 $X=613800 $Y=1722718
X45 1003 3 1034 955 1 NOR2BX1 $T=561660 1672720 1 0 $X=561658 $Y=1667280
X46 33 1121 1110 1098 3 1 1064 ADDFX2 $T=595980 1733200 0 180 $X=582120 $Y=1727760
X47 1284 39 1227 1121 3 1 1219 ADDFX2 $T=630960 1763440 0 180 $X=617100 $Y=1758000
X48 1228 1249 1245 36 3 1 1175 ADDFX2 $T=634920 1642480 1 180 $X=621060 $Y=1642078
X49 1262 1255 38 37 3 1 1228 ADDFX2 $T=635580 1622320 0 180 $X=621720 $Y=1616880
X50 44 42 41 40 3 1 1262 ADDFX2 $T=650100 1632400 0 180 $X=636240 $Y=1626960
X51 1304 47 1283 1277 3 1 1191 ADDFX2 $T=652740 1733200 1 180 $X=638880 $Y=1732798
X52 1281 50 1277 1280 3 1 1174 ADDFX2 $T=654060 1702960 0 180 $X=640200 $Y=1697520
X53 41 52 1291 1281 3 1 1205 ADDFX2 $T=654720 1702960 1 180 $X=640860 $Y=1702558
X54 1292 1287 1286 1282 3 1 1204 ADDFX2 $T=655380 1682800 1 180 $X=641520 $Y=1682398
X55 52 53 45 1290 3 1 1286 ADDFX2 $T=657360 1662640 0 180 $X=643500 $Y=1657200
X56 43 54 46 1292 3 1 1283 ADDFX2 $T=657360 1723120 1 180 $X=643500 $Y=1722718
X57 63 53 48 1190 3 1 1227 ADDFX2 $T=657360 1743280 0 180 $X=643500 $Y=1737840
X58 42 54 45 1304 3 1 1284 ADDFX2 $T=658680 1763440 0 180 $X=644820 $Y=1758000
X59 1329 1290 1326 1245 3 1 1279 ADDFX2 $T=660000 1642480 0 180 $X=646140 $Y=1637040
X60 75 46 61 1249 3 1 1326 ADDFX2 $T=665280 1652560 0 180 $X=651420 $Y=1647120
X61 51 1291 44 3 1 1287 ADDHXL $T=652740 1713040 1 180 $X=645480 $Y=1712638
X62 3 1001 957 954 1 NOR2XL $T=551100 1713040 0 180 $X=549120 $Y=1707600
X63 16 954 924 1 923 3 OAI2BB1X1 $T=538560 1713040 0 180 $X=535260 $Y=1707600
X64 938 922 941 1 956 3 OAI2BB1X1 $T=540540 1662640 0 0 $X=540538 $Y=1662238
X65 938 1005 1006 1 1048 3 OAI2BB1X1 $T=553080 1662640 0 0 $X=553078 $Y=1662238
X66 20 16 25 1 32 3 OAI2BB1X1 $T=569580 1773520 0 0 $X=569578 $Y=1773118
X67 30 1093 1049 1 1044 3 OAI2BB1X1 $T=583440 1773520 0 180 $X=580140 $Y=1768080
X68 939 1 937 3 908 NAND2BXL $T=540540 1702960 1 180 $X=537900 $Y=1702558
X69 1001 1 1033 3 1017 NAND2BXL $T=561660 1713040 1 180 $X=559020 $Y=1712638
X70 1034 1 1062 3 1050 NAND2BXL $T=571560 1662640 0 180 $X=568920 $Y=1657200
X71 1101 1 1095 3 1080 NAND2BXL $T=584100 1642480 1 180 $X=581460 $Y=1642078
X72 16 938 1 3 CLKBUFX3 $T=540540 1713040 1 0 $X=540538 $Y=1707600
X73 1001 1007 1067 1064 3 1 924 AOI2BB2X1 $T=574200 1723120 0 180 $X=569580 $Y=1717680
X74 1204 1187 1174 1122 3 1 1120 ADDFHX1 $T=613800 1692880 1 180 $X=598620 $Y=1692478
X75 1219 35 34 1067 3 1 1079 ADDFHX1 $T=627000 1773520 0 180 $X=611820 $Y=1768080
X76 1282 1280 1279 1129 3 1 1173 ADDFHX1 $T=655380 1672720 0 180 $X=640200 $Y=1667280
X77 1189 1 1188 3 1192 1187 NAND3X1 $T=606540 1713040 0 180 $X=603900 $Y=1707600
X78 43 45 54 1255 1 3 1329 CMPR32X1 $T=646140 1622320 1 0 $X=646138 $Y=1616880
.ENDS
***************************************
.SUBCKT OAI2BB2X2 A0N A1N Y B0 B1 VSS VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB1X2 A0N A1N Y VSS B0 VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDFHX2 A B CI CO VDD VSS S
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDFHX4 A B CI CO S VSS VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_76 1 3 22 23 24 25 26 27 28 29 30 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 55 56 57 58 59 60 61
+ 70 71 72 73 74 75 76 77 86 88 89 345 346
** N=4604 EP=53 IP=428 FDC=0
X0 1186 3 1169 1 1164 NAND2X1 $T=565620 1854160 0 180 $X=563640 $Y=1848720
X1 26 3 1202 1 1168 NAND2X1 $T=572220 1793680 1 0 $X=572218 $Y=1788240
X2 1238 3 1224 1 1254 NAND2X1 $T=585420 1803760 1 0 $X=585418 $Y=1798320
X3 1339 3 1343 1 1341 NAND2X1 $T=609840 1894480 1 180 $X=607860 $Y=1894078
X4 1375 3 1339 1 1338 NAND2X1 $T=616440 1874320 1 180 $X=614460 $Y=1873918
X5 1164 3 1 1071 INVX1 $T=550440 1813840 0 180 $X=549120 $Y=1808400
X6 28 3 1 1202 INVX1 $T=583440 1793680 1 0 $X=583438 $Y=1788240
X7 1254 3 1 29 INVX1 $T=584760 1783600 0 180 $X=583440 $Y=1778160
X8 1 1185 1166 1167 3 NOR2X1 $T=562980 1844080 0 180 $X=561000 $Y=1838640
X9 1 1167 1088 26 3 NOR2X1 $T=563640 1823920 1 180 $X=561660 $Y=1823518
X10 1 1238 1224 28 3 NOR2X1 $T=580140 1803760 0 180 $X=578160 $Y=1798320
X11 1169 1186 3 1 1088 NOR2X2 $T=566940 1864240 0 180 $X=563640 $Y=1858800
X12 1202 1 1254 3 1270 AND2X2 $T=595320 1783600 0 0 $X=595318 $Y=1783198
X13 1088 1071 3 1 1070 OR2X2 $T=545820 1813840 0 180 $X=543180 $Y=1808400
X14 1375 3 1 1343 1340 NAND2XL $T=608520 1874320 1 180 $X=606540 $Y=1873918
X15 42 3 1 41 1453 NAND2XL $T=636900 1975120 0 180 $X=634920 $Y=1969680
X16 48 3 1 41 1456 NAND2XL $T=636900 1985200 1 180 $X=634920 $Y=1984798
X17 39 3 1 41 1553 NAND2XL $T=652740 1985200 0 180 $X=650760 $Y=1979760
X18 70 3 1 45 61 NAND2XL $T=655380 1924720 0 180 $X=653400 $Y=1919280
X19 41 3 1 49 1550 NAND2XL $T=660660 1975120 0 180 $X=658680 $Y=1969680
X20 1168 22 3 1184 1 25 OAI21X2 $T=561660 1783600 0 0 $X=561658 $Y=1783198
X21 1088 3 22 1164 1 1203 OAI21X4 $T=560340 1813840 1 0 $X=560338 $Y=1808400
X22 1070 22 1 3 23 XOR2X2 $T=554400 1803760 1 0 $X=554398 $Y=1798320
X23 1270 32 1 3 33 XOR2X2 $T=593340 1783600 1 0 $X=593338 $Y=1778160
X24 1219 1203 1 3 30 XNOR2X2 $T=574860 1813840 1 0 $X=574858 $Y=1808400
X25 1448 39 3 1 1451 XOR2X1 $T=630960 1965040 0 0 $X=630958 $Y=1964638
X26 49 41 3 1 1448 XOR2X1 $T=648120 1965040 0 180 $X=642840 $Y=1959600
X27 71 45 3 1 88 XOR2X1 $T=656040 1944880 0 0 $X=656038 $Y=1944478
X28 88 70 3 1 1482 XOR2X1 $T=662640 1934800 1 180 $X=657360 $Y=1934398
X29 1412 1398 1379 34 1 3 1224 ADDFX2 $T=621060 1803760 0 180 $X=607200 $Y=1798320
X30 1489 36 1417 35 1 3 1379 ADDFX2 $T=633600 1823920 0 180 $X=619740 $Y=1818480
X31 1551 1451 37 1434 1 3 1339 ADDFX2 $T=638880 1904560 0 180 $X=625020 $Y=1899120
X32 46 1452 38 1436 1 3 1343 ADDFX2 $T=639540 1934800 0 180 $X=625680 $Y=1929360
X33 1482 1455 1436 1412 1 3 1418 ADDFX2 $T=640200 1904560 1 180 $X=626340 $Y=1904158
X34 1552 51 44 1375 1 3 1472 ADDFX2 $T=652080 1874320 0 180 $X=638220 $Y=1868880
X35 59 1508 1486 1417 1 3 1473 ADDFX2 $T=652740 1834000 1 180 $X=638880 $Y=1833598
X36 45 50 39 1556 1 3 1507 ADDFX2 $T=643500 1793680 1 0 $X=643498 $Y=1788240
X37 52 1556 1490 47 1 3 43 ADDFX2 $T=657360 1783600 0 180 $X=643500 $Y=1778160
X38 74 1491 1507 1490 1 3 1398 ADDFX2 $T=657360 1793680 1 180 $X=643500 $Y=1793278
X39 76 60 48 1491 1 3 1486 ADDFX2 $T=657360 1803760 1 180 $X=643500 $Y=1803358
X40 72 49 55 52 1 3 1489 ADDFX2 $T=660000 1823920 0 180 $X=646140 $Y=1818480
X41 56 1557 77 37 1 3 89 ADDFX2 $T=650760 1894480 0 0 $X=650758 $Y=1894078
X42 45 71 86 38 1 3 77 ADDFX2 $T=651420 1934800 1 0 $X=651418 $Y=1929360
X43 49 42 72 1557 1 3 57 ADDFX2 $T=665280 1894480 0 180 $X=651420 $Y=1889040
X44 76 72 73 1455 1 3 1551 ADDFX2 $T=665280 1904560 1 180 $X=651420 $Y=1904158
X45 1185 1166 3 1 1219 XNOR2X1 $T=581460 1834000 1 180 $X=576180 $Y=1833598
X46 1375 1343 1339 3 1 1169 XOR3X2 $T=610500 1884400 1 180 $X=598620 $Y=1883998
X47 42 41 48 3 1 1552 XOR3X2 $T=636900 1934800 0 0 $X=636898 $Y=1934398
X48 1340 3 1338 1 1341 1185 NAND3X1 $T=601260 1874320 1 180 $X=598620 $Y=1873918
X49 1453 3 40 1 1456 1452 NAND3X1 $T=634920 1985200 1 0 $X=634918 $Y=1979760
X50 58 3 1553 1 1550 1508 NAND3X1 $T=652080 1975120 0 180 $X=649440 $Y=1969680
X51 1166 1185 24 1167 1164 3 1 OAI2BB2X2 $T=567600 1834000 1 180 $X=561000 $Y=1833598
X52 28 27 1184 3 29 1 AOI2BB1X2 $T=574860 1783600 1 0 $X=574858 $Y=1778160
X53 1473 1434 1418 1238 1 3 1166 ADDFHX2 $T=644160 1854160 0 180 $X=621720 $Y=1848720
X54 89 75 1472 1186 53 3 1 ADDFHX4 $T=671220 1864240 1 180 $X=648120 $Y=1863838
.ENDS
***************************************
.SUBCKT ICV_75 2 4 39 40 41 303 304
** N=5170 EP=7 IP=7 FDC=0
X0 41 2 4 40 39 NAND2XL $T=638220 1995280 1 180 $X=636240 $Y=1994878
.ENDS
***************************************
.SUBCKT ICV_74
** N=3894 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_73
** N=3777 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_72
** N=5059 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_71
** N=3424 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_70
** N=4125 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_69 3 4 5 6 7 8
** N=17 EP=6 IP=12 FDC=0
X0 3 5 PDIDGZ $T=504100 3289640 0 180 $X=476420 $Y=3104640
X1 4 6 PDIDGZ $T=663650 3289640 0 180 $X=635970 $Y=3104640
.ENDS
***************************************
.SUBCKT OR2X1 A B VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX3 A VDD Y VSS
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2X1 A B VDD VSS Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB1X4 A0N A1N B0 VDD Y VSS
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22X1 B1 B0 VDD A0 A1 Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB2X1 A0N A1N B1 B0 VSS VDD Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDFXL B A CI CO VSS VDD S
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2XL B A VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2X4 A B Y VDD VSS
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB1X4 A1N A0N B0 VSS VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX8 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MX2X4 B S0 A Y VDD VSS
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB2X4 A1N A0N B1 VSS B0 Y VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2BX2 AN B Y VSS VDD
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB1X2 A1N A0N B0 Y VDD VSS
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND3X1 A B C VSS VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND3X2 A B C VSS VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3BXL AN VSS C B VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2BX2 AN B Y VSS VDD
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2XL B A VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3X2 VDD A Y B C VSS
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRHQXL CK SE SI D RN VDD VSS Q
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX3 A VDD Y VSS
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI221X1 B1 B0 A0 VDD A1 VSS C0 Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI32XL A2 A1 A0 VDD B0 B1 VSS Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX4 A Y VDD VSS
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI222X2 C0 C1 VDD B1 B0 A0 A1 Y VSS
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22X1 B1 B0 VSS A0 A1 VDD Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2BXL AN VDD B Y VSS
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR3BX1 AN VDD C B VSS Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI211X1 A1 VDD A0 C0 VSS B0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI32X1 A2 A1 A0 VSS B0 B1 VDD Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB1X1 A0N A1N VSS VDD B0 Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI222X1 C0 C1 VDD B1 B0 A0 Y A1 VSS
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI2X1 S0 B Y A VSS VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI211X1 A1 A0 VSS C0 VDD B0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNOR3X2 A B C VSS VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22XL B1 VDD B0 A0 A1 Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB1XL A0N A1N VSS B0 VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI211X2 A1 A0 VDD B0 VSS C0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI211X2 A1 A0 VSS VDD B0 C0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4BX1 AN VDD D C B Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI31X4 A2 A1 A0 B0 VDD VSS Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX4 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR4X2 A B C VSS D VDD Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2BX4 AN B VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDHX4 B S A CO VDD VSS
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI32X1 A2 A1 A0 VDD B0 B1 VSS Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI33X1 B2 B1 VSS B0 A0 A1 A2 VDD Y
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3XL A B C VDD VSS Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22XL B1 B0 VSS A0 A1 Y VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI31X1 A2 A1 A0 VSS B0 VDD Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND3X4 A B C Y VSS VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4X1 VDD D C B A Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3XL C VSS B VDD A Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI221XL B1 B0 VDD A0 A1 VSS C0 Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB1XL A1N A0N B0 VSS Y VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222X1 B1 B0 VSS A0 A1 VDD C1 C0 Y
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX8 A VSS Y VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR3X1 C VDD B VSS A Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI222X4 C1 C0 B1 B0 A0 A1 Y VSS VDD
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRXL CK SE SI D RN QN VSS VDD Q
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2BX4 AN B VDD VSS Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4X2 A VSS B C D Y VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4XL D VDD C B A Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4BBX2 AN D C BN VSS Y VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3BX2 Y B C VDD VSS AN
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222XL B1 B0 A0 VSS A1 VDD C1 C0 Y
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2X4 A B VSS VDD Y
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MX2X1 S0 B A VSS VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX12 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX8 A VDD VSS Y
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22X2 B0 B1 VDD A0 A1 Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX16 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI2X4 A Y S0 B VSS VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_62 1 3 42 45 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68
+ 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128
+ 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188
+ 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208
+ 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228
+ 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248
+ 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263 264 265 266 267 268
+ 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286 287 288
+ 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304 305 306 307 308
+ 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 326 327 328
+ 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347 348
+ 349 350 351 352 353 354 355 356 357 360 361 362 363 364 365 366 367 368 369 370
+ 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390
+ 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410
+ 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430
+ 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 499 500 501 502 503 504 505 506 507 508 509 510 511
+ 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 529 530 531 532
+ 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552
+ 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572
+ 573 574 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591 592
+ 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610 611 612
+ 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629 630 631 632
+ 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648 649 650 651 652
+ 653 654 655 656 657 658 659 660 661 662 663 664 666 667 668 669 670 671 672 673
+ 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690 691 692 693
+ 694 695 696 697 1480 1481
** N=46430 EP=646 IP=17378 FDC=0
X0 67 1 1511 3 1543 NAND2X1 $T=671220 1269520 1 180 $X=669240 $Y=1269118
X1 64 1 1541 3 1576 NAND2X1 $T=673200 1219120 1 0 $X=673198 $Y=1213680
X2 1597 1 1549 3 1545 NAND2X1 $T=676500 1279600 0 180 $X=674520 $Y=1274160
X3 1567 1 1508 3 1745 NAND2X1 $T=679800 1309840 0 0 $X=679798 $Y=1309438
X4 1602 1 1606 3 1609 NAND2X1 $T=682440 1259440 1 0 $X=682438 $Y=1254000
X5 1611 1 1608 3 1607 NAND2X1 $T=684420 1380400 0 180 $X=682440 $Y=1374960
X6 68 1 1601 3 1603 NAND2X1 $T=689040 1229200 0 0 $X=689038 $Y=1228798
X7 1636 1 1634 3 1631 NAND2X1 $T=691020 1350160 1 180 $X=689040 $Y=1349758
X8 1669 1 72 3 1608 NAND2X1 $T=695640 1380400 1 180 $X=693660 $Y=1379998
X9 1660 1 72 3 1634 NAND2X1 $T=695640 1370320 0 0 $X=695638 $Y=1369918
X10 1549 1 1602 3 1748 NAND2X1 $T=701580 1249360 1 0 $X=701578 $Y=1243920
X11 1887 1 1750 3 1746 NAND2X1 $T=712800 1380400 1 180 $X=710820 $Y=1379998
X12 1808 1 1814 3 1780 NAND2X1 $T=713460 1249360 1 0 $X=713458 $Y=1243920
X13 1870 1 1602 3 1840 NAND2X1 $T=720060 1249360 1 180 $X=718080 $Y=1248958
X14 1846 1 1847 3 1744 NAND2X1 $T=719400 1269520 1 0 $X=719398 $Y=1264080
X15 81 1 1897 3 1846 NAND2X1 $T=726000 1279600 1 0 $X=725998 $Y=1274160
X16 79 1 1865 3 1915 NAND2X1 $T=727980 1289680 1 180 $X=726000 $Y=1289278
X17 1915 1 1870 3 1981 NAND2X1 $T=729300 1249360 0 0 $X=729298 $Y=1248958
X18 1846 1 1942 3 1914 NAND2X1 $T=731940 1269520 1 0 $X=731938 $Y=1264080
X19 2012 1 83 3 1898 NAND2X1 $T=737880 1400560 1 180 $X=735900 $Y=1400158
X20 1927 1 1985 3 85 NAND2X1 $T=738540 1168720 1 0 $X=738538 $Y=1163280
X21 1980 1 1887 3 1924 NAND2X1 $T=738540 1380400 0 0 $X=738538 $Y=1379998
X22 2108 1 1782 3 1956 NAND2X1 $T=744480 1360240 0 180 $X=742500 $Y=1354800
X23 88 1 86 3 1917 NAND2X1 $T=757020 1430800 1 0 $X=757018 $Y=1425360
X24 89 1 2182 3 1989 NAND2X1 $T=766920 1420720 0 0 $X=766918 $Y=1420318
X25 2245 1 2208 3 1980 NAND2X1 $T=768900 1390480 1 180 $X=766920 $Y=1390078
X26 2241 1 2212 3 2170 NAND2X1 $T=770220 1219120 0 180 $X=768240 $Y=1213680
X27 2236 1 2232 3 2145 NAND2X1 $T=771540 1330000 1 180 $X=769560 $Y=1329598
X28 2275 1 2241 3 2179 NAND2X1 $T=774180 1239280 0 180 $X=772200 $Y=1233840
X29 91 1 2269 3 2202 NAND2X1 $T=776160 1168720 1 0 $X=776158 $Y=1163280
X30 2305 1 2241 3 2302 NAND2X1 $T=780780 1209040 1 180 $X=778800 $Y=1208638
X31 2307 1 2282 3 2167 NAND2X1 $T=782100 1370320 0 0 $X=782098 $Y=1369918
X32 2309 1 2242 3 2235 NAND2X1 $T=782760 1299760 0 0 $X=782758 $Y=1299358
X33 2374 1 2370 3 2275 NAND2X1 $T=792660 1239280 1 180 $X=790680 $Y=1238878
X34 2404 1 2371 3 2285 NAND2X1 $T=798600 1279600 0 0 $X=798598 $Y=1279198
X35 2543 1 2518 3 2346 NAND2X1 $T=818400 1279600 1 0 $X=818398 $Y=1274160
X36 2171 1 2619 3 2642 NAND2X1 $T=832920 1178800 1 0 $X=832918 $Y=1173360
X37 2642 1 2635 3 2764 NAND2X1 $T=838860 1178800 1 0 $X=838858 $Y=1173360
X38 2140 1 2671 3 2672 NAND2X1 $T=844140 1198960 0 0 $X=844138 $Y=1198558
X39 115 1 2869 3 2842 NAND2X1 $T=871860 1209040 1 0 $X=871858 $Y=1203600
X40 2922 1 2937 3 3008 NAND2X1 $T=885060 1249360 0 0 $X=885058 $Y=1248958
X41 54 1 2949 3 3062 NAND2X1 $T=887700 1390480 0 0 $X=887698 $Y=1390078
X42 3162 1 3137 3 121 NAND2X1 $T=919380 1158640 1 180 $X=917400 $Y=1158238
X43 3214 1 3162 3 3092 NAND2X1 $T=932580 1178800 0 180 $X=930600 $Y=1173360
X44 126 1 3349 3 3197 NAND2X1 $T=954360 1158640 1 0 $X=954358 $Y=1153200
X45 3403 1 3358 3 3356 NAND2X1 $T=956340 1299760 0 180 $X=954360 $Y=1294320
X46 3445 1 3408 3 3372 NAND2X1 $T=962940 1410640 1 180 $X=960960 $Y=1410238
X47 141 1 140 3 3414 NAND2X1 $T=975480 1229200 0 0 $X=975478 $Y=1228798
X48 3550 1 3505 3 3445 NAND2X1 $T=980760 1410640 1 180 $X=978780 $Y=1410238
X49 137 1 3534 3 3435 NAND2X1 $T=985380 1360240 1 0 $X=985378 $Y=1354800
X50 145 1 144 3 3465 NAND2X1 $T=987360 1299760 0 180 $X=985380 $Y=1294320
X51 146 1 3557 3 3437 NAND2X1 $T=990000 1309840 0 180 $X=988020 $Y=1304400
X52 148 1 149 3 3478 NAND2X1 $T=995280 1309840 0 0 $X=995278 $Y=1309438
X53 3588 1 3672 3 3712 NAND2X1 $T=1002540 1340080 0 0 $X=1002538 $Y=1339678
X54 3713 1 3733 3 3557 NAND2X1 $T=1008480 1400560 0 0 $X=1008478 $Y=1400158
X55 3731 1 158 3 3733 NAND2X1 $T=1010460 1410640 1 0 $X=1010458 $Y=1405200
X56 3739 1 3670 3 161 NAND2X1 $T=1012440 1148560 0 180 $X=1010460 $Y=1143120
X57 3854 1 3732 3 3794 NAND2X1 $T=1019040 1279600 1 180 $X=1017060 $Y=1279198
X58 3841 1 3796 3 3615 NAND2X1 $T=1023000 1188880 0 180 $X=1021020 $Y=1183440
X59 3857 1 3856 3 3855 NAND2X1 $T=1032240 1370320 0 180 $X=1030260 $Y=1364880
X60 3801 1 3854 3 3741 NAND2X1 $T=1030920 1279600 0 0 $X=1030918 $Y=1279198
X61 3877 1 3906 3 3699 NAND2X1 $T=1034880 1330000 0 0 $X=1034878 $Y=1329598
X62 3902 1 3875 3 3698 NAND2X1 $T=1038180 1249360 1 0 $X=1038178 $Y=1243920
X63 3898 1 3856 3 3867 NAND2X1 $T=1038840 1370320 0 0 $X=1038838 $Y=1369918
X64 3922 1 3905 3 3866 NAND2X1 $T=1041480 1229200 1 180 $X=1039500 $Y=1228798
X65 3921 1 3904 3 3711 NAND2X1 $T=1040820 1168720 1 0 $X=1040818 $Y=1163280
X66 4021 1 3951 3 3898 NAND2X1 $T=1047420 1360240 0 180 $X=1045440 $Y=1354800
X67 3955 1 3857 3 3834 NAND2X1 $T=1048080 1370320 0 0 $X=1048078 $Y=1369918
X68 4022 1 3957 3 3836 NAND2X1 $T=1050720 1319920 0 0 $X=1050718 $Y=1319518
X69 4031 1 3903 3 3804 NAND2X1 $T=1054020 1259440 0 0 $X=1054018 $Y=1259038
X70 4026 1 4060 3 4057 NAND2X1 $T=1060620 1168720 1 180 $X=1058640 $Y=1168318
X71 4026 1 4086 3 4030 NAND2X1 $T=1059960 1178800 1 0 $X=1059958 $Y=1173360
X72 4089 1 4093 3 3955 NAND2X1 $T=1064580 1370320 0 0 $X=1064578 $Y=1369918
X73 4266 1 4146 3 4090 NAND2X1 $T=1072500 1390480 1 180 $X=1070520 $Y=1390078
X74 4141 1 4149 3 4152 NAND2X1 $T=1071840 1279600 1 0 $X=1071838 $Y=1274160
X75 4215 1 4186 3 175 NAND2X1 $T=1080420 1420720 0 180 $X=1078440 $Y=1415280
X76 4141 1 4209 3 4156 NAND2X1 $T=1090320 1279600 1 0 $X=1090318 $Y=1274160
X77 4410 1 4367 3 4411 NAND2X1 $T=1116060 1319920 1 180 $X=1114080 $Y=1319518
X78 211 1 4507 3 4524 NAND2X1 $T=1141800 1420720 0 180 $X=1139820 $Y=1415280
X79 4410 1 4460 3 4455 NAND2X1 $T=1145100 1319920 0 0 $X=1145098 $Y=1319518
X80 192 1 217 3 4674 NAND2X1 $T=1165560 1420720 1 180 $X=1163580 $Y=1420318
X81 4459 1 191 3 4669 NAND2X1 $T=1179420 1209040 0 0 $X=1179418 $Y=1208638
X82 199 1 230 3 5019 NAND2X1 $T=1217700 1229200 1 180 $X=1215720 $Y=1228798
X83 247 1 187 3 5226 NAND2X1 $T=1236840 1198960 0 0 $X=1236838 $Y=1198558
X84 5191 1 5463 3 5459 NAND2X1 $T=1270500 1198960 0 0 $X=1270498 $Y=1198558
X85 5835 1 288 3 5832 NAND2X1 $T=1345740 1229200 1 180 $X=1343760 $Y=1228798
X86 290 1 5835 3 5842 NAND2X1 $T=1345740 1239280 0 180 $X=1343760 $Y=1233840
X87 290 1 288 3 5839 NAND2X1 $T=1347060 1259440 0 180 $X=1345080 $Y=1254000
X88 284 1 288 3 5925 NAND2X1 $T=1354320 1350160 1 0 $X=1354318 $Y=1344720
X89 5997 1 6000 3 6007 NAND2X1 $T=1367520 1330000 1 0 $X=1367518 $Y=1324560
X90 6007 1 6088 3 6104 NAND2X1 $T=1380720 1330000 1 0 $X=1380718 $Y=1324560
X91 6068 1 6039 3 6192 NAND2X1 $T=1383360 1319920 1 0 $X=1383358 $Y=1314480
X92 6044 1 6253 3 6281 NAND2X1 $T=1401180 1239280 1 0 $X=1401178 $Y=1233840
X93 5614 1 6087 3 6279 NAND2X1 $T=1401180 1289680 1 0 $X=1401178 $Y=1284240
X94 6165 1 6277 3 6278 NAND2X1 $T=1405140 1198960 1 0 $X=1405138 $Y=1193520
X95 6192 1 6095 3 6283 NAND2X1 $T=1409100 1319920 1 0 $X=1409098 $Y=1314480
X96 6149 1 6251 3 6306 NAND2X1 $T=1410420 1229200 1 0 $X=1410418 $Y=1223760
X97 307 1 3379 3 6379 NAND2X1 $T=1414380 1410640 1 180 $X=1412400 $Y=1410238
X98 6160 1 6335 3 6368 NAND2X1 $T=1415700 1168720 0 0 $X=1415698 $Y=1168318
X99 6440 1 5948 3 308 NAND2X1 $T=1419000 1420720 1 180 $X=1417020 $Y=1420318
X100 6422 1 6405 3 6429 NAND2X1 $T=1430880 1198960 1 0 $X=1430878 $Y=1193520
X101 5711 1 6378 3 6433 NAND2X1 $T=1432860 1279600 0 0 $X=1432858 $Y=1279198
X102 6368 1 6405 3 6567 NAND2X1 $T=1435500 1168720 0 0 $X=1435498 $Y=1168318
X103 6278 1 6422 3 6569 NAND2X1 $T=1443420 1198960 1 0 $X=1443418 $Y=1193520
X104 6422 1 6505 3 6591 NAND2X1 $T=1446060 1188880 0 0 $X=1446058 $Y=1188478
X105 6593 1 6572 3 6640 NAND2X1 $T=1457280 1350160 0 0 $X=1457278 $Y=1349758
X106 5649 1 6595 3 6660 NAND2X1 $T=1457940 1259440 0 0 $X=1457938 $Y=1259038
X107 6434 1 6597 3 6659 NAND2X1 $T=1464540 1400560 1 0 $X=1464538 $Y=1395120
X108 6005 1 6627 3 6735 NAND2X1 $T=1469160 1209040 0 0 $X=1469158 $Y=1208638
X109 321 1 3359 3 6763 NAND2X1 $T=1471140 1330000 1 180 $X=1469160 $Y=1329598
X110 6693 1 6695 3 6752 NAND2X1 $T=1470480 1158640 1 0 $X=1470478 $Y=1153200
X111 6696 1 3274 3 6732 NAND2X1 $T=1474440 1269520 1 180 $X=1472460 $Y=1269118
X112 6798 1 6759 3 6803 NAND2X1 $T=1489620 1340080 1 0 $X=1489618 $Y=1334640
X113 322 1 3352 3 6940 NAND2X1 $T=1492920 1340080 0 0 $X=1492918 $Y=1339678
X114 293 1 327 3 330 NAND2X1 $T=1503480 1138480 0 0 $X=1503478 $Y=1138078
X115 6702 1 6737 3 6952 NAND2X1 $T=1505460 1158640 1 0 $X=1505458 $Y=1153200
X116 6941 1 6948 3 6944 NAND2X1 $T=1508100 1390480 0 0 $X=1508098 $Y=1390078
X117 6979 1 6978 3 7058 NAND2X1 $T=1517340 1209040 0 0 $X=1517338 $Y=1208638
X118 7000 1 3013 3 7028 NAND2X1 $T=1518000 1229200 1 0 $X=1517998 $Y=1223760
X119 6978 1 7028 3 7030 NAND2X1 $T=1523280 1219120 0 0 $X=1523278 $Y=1218718
X120 6839 1 7095 3 7074 NAND2X1 $T=1529880 1350160 0 0 $X=1529878 $Y=1349758
X121 6725 1 7162 3 7056 NAND2X1 $T=1542420 1410640 1 0 $X=1542418 $Y=1405200
X122 7292 1 7103 3 7321 NAND2X1 $T=1560240 1360240 0 180 $X=1558260 $Y=1354800
X123 7180 1 7393 3 7286 NAND2X1 $T=1576740 1330000 0 0 $X=1576738 $Y=1329598
X124 7415 1 7406 3 7384 NAND2X1 $T=1580040 1239280 1 180 $X=1578060 $Y=1238878
X125 6922 1 7389 3 7471 NAND2X1 $T=1582020 1299760 0 0 $X=1582018 $Y=1299358
X126 7478 1 7071 3 7418 NAND2X1 $T=1591920 1198960 0 0 $X=1591918 $Y=1198558
X127 7502 1 7177 3 7543 NAND2X1 $T=1600500 1319920 0 0 $X=1600498 $Y=1319518
X128 7771 1 7754 3 6100 NAND2X1 $T=1633500 1390480 0 180 $X=1631520 $Y=1385040
X129 7806 1 7655 3 7765 NAND2X1 $T=1637460 1198960 1 180 $X=1635480 $Y=1198558
X130 7760 1 7288 3 7797 NAND2X1 $T=1639440 1229200 1 0 $X=1639438 $Y=1223760
X131 7930 1 7795 3 6370 NAND2X1 $T=1641420 1370320 0 180 $X=1639440 $Y=1364880
X132 7527 1 7833 3 7953 NAND2X1 $T=1646700 1259440 0 180 $X=1644720 $Y=1254000
X133 7924 1 7802 3 7928 NAND2X1 $T=1654620 1259440 1 180 $X=1652640 $Y=1259038
X134 7951 1 361 3 7922 NAND2X1 $T=1654620 1400560 1 180 $X=1652640 $Y=1400158
X135 7987 1 8035 3 8045 NAND2X1 $T=1671120 1198960 0 0 $X=1671118 $Y=1198558
X136 7479 1 8036 3 7950 NAND2X1 $T=1671120 1259440 1 0 $X=1671118 $Y=1254000
X137 7527 1 7962 3 8126 NAND2X1 $T=1679700 1239280 1 0 $X=1679698 $Y=1233840
X138 7527 1 8098 3 8362 NAND2X1 $T=1683660 1229200 0 0 $X=1683658 $Y=1228798
X139 8152 1 6342 3 8100 NAND2X1 $T=1686960 1360240 0 180 $X=1684980 $Y=1354800
X140 8168 1 6671 3 8243 NAND2X1 $T=1694880 1309840 1 180 $X=1692900 $Y=1309438
X141 8149 1 8274 3 385 NAND2X1 $T=1709400 1138480 1 180 $X=1707420 $Y=1138078
X142 8149 1 8296 3 8309 NAND2X1 $T=1711380 1158640 1 0 $X=1711378 $Y=1153200
X143 8340 1 8338 3 6371 NAND2X1 $T=1719960 1340080 1 180 $X=1717980 $Y=1339678
X144 8149 1 8304 3 8415 NAND2X1 $T=1725240 1239280 1 0 $X=1725238 $Y=1233840
X145 8413 1 8381 3 6106 NAND2X1 $T=1727880 1330000 1 180 $X=1725900 $Y=1329598
X146 8149 1 8400 3 398 NAND2X1 $T=1728540 1138480 0 0 $X=1728538 $Y=1138078
X147 8303 1 387 3 8310 NAND2X1 $T=1728540 1148560 0 0 $X=1728538 $Y=1148158
X148 8311 1 387 3 8402 NAND2X1 $T=1728540 1239280 1 0 $X=1728538 $Y=1233840
X149 8574 1 6568 3 8477 NAND2X1 $T=1753620 1289680 0 180 $X=1751640 $Y=1284240
X150 8627 1 7010 3 8633 NAND2X1 $T=1758900 1209040 1 180 $X=1756920 $Y=1208638
X151 8628 1 6852 3 8622 NAND2X1 $T=1764840 1269520 1 0 $X=1764838 $Y=1264080
X152 8656 1 7352 3 8658 NAND2X1 $T=1769460 1188880 1 180 $X=1767480 $Y=1188478
X153 8863 1 6825 3 8729 NAND2X1 $T=1799820 1249360 0 180 $X=1797840 $Y=1243920
X154 448 1 447 3 8916 NAND2X1 $T=1809720 1340080 0 180 $X=1807740 $Y=1334640
X155 8919 1 7264 3 8862 NAND2X1 $T=1812360 1138480 0 0 $X=1812358 $Y=1138078
X156 8619 1 8975 3 8977 NAND2X1 $T=1820280 1319920 1 0 $X=1820278 $Y=1314480
X157 8433 1 9043 3 8984 NAND2X1 $T=1823580 1299760 0 0 $X=1823578 $Y=1299358
X158 456 1 455 3 8981 NAND2X1 $T=1829520 1390480 1 180 $X=1827540 $Y=1390078
X159 8649 1 9038 3 9130 NAND2X1 $T=1831500 1340080 1 0 $X=1831498 $Y=1334640
X160 8591 1 9062 3 9058 NAND2X1 $T=1834800 1350160 1 0 $X=1834798 $Y=1344720
X161 8625 1 9068 3 9076 NAND2X1 $T=1838100 1330000 1 0 $X=1838098 $Y=1324560
X162 474 1 473 3 9190 NAND2X1 $T=1858560 1138480 1 180 $X=1856580 $Y=1138078
X163 8596 1 9236 3 9207 NAND2X1 $T=1861860 1259440 1 0 $X=1861858 $Y=1254000
X164 8679 1 9286 3 9343 NAND2X1 $T=1869780 1239280 0 0 $X=1869778 $Y=1238878
X165 8620 1 9297 3 9327 NAND2X1 $T=1871100 1259440 1 0 $X=1871098 $Y=1254000
X166 9326 1 9324 3 478 NAND2X1 $T=1879680 1269520 1 180 $X=1877700 $Y=1269118
X167 484 1 481 3 480 NAND2X1 $T=1881000 1138480 1 180 $X=1879020 $Y=1138078
X168 8414 1 9405 3 9404 NAND2X1 $T=1890900 1209040 1 0 $X=1890898 $Y=1203600
X169 485 1 486 3 9383 NAND2X1 $T=1894200 1400560 0 0 $X=1894198 $Y=1400158
X170 9437 1 9444 3 489 NAND2X1 $T=1898160 1259440 0 0 $X=1898158 $Y=1259038
X171 435 1 9507 3 9529 NAND2X1 $T=1898160 1289680 1 0 $X=1898158 $Y=1284240
X172 492 1 491 3 9438 NAND2X1 $T=1902120 1370320 0 180 $X=1900140 $Y=1364880
X173 9504 1 493 3 9567 NAND2X1 $T=1903440 1209040 0 0 $X=1903438 $Y=1208638
X174 9443 1 493 3 9565 NAND2X1 $T=1904760 1188880 0 0 $X=1904758 $Y=1188478
X175 431 1 493 3 9533 NAND2X1 $T=1908720 1299760 1 0 $X=1908718 $Y=1294320
X176 435 1 9572 3 9593 NAND2X1 $T=1915980 1209040 1 180 $X=1914000 $Y=1208638
X177 435 1 9595 3 9573 NAND2X1 $T=1919280 1188880 0 0 $X=1919278 $Y=1188478
X178 9328 1 493 3 9621 NAND2X1 $T=1919280 1289680 0 0 $X=1919278 $Y=1289278
X179 449 1 9592 3 9623 NAND2X1 $T=1921920 1319920 0 180 $X=1919940 $Y=1314480
X180 9623 1 9631 3 9634 NAND2X1 $T=1921920 1219120 1 0 $X=1921918 $Y=1213680
X181 449 1 9664 3 9570 NAND2X1 $T=1927860 1309840 1 0 $X=1927858 $Y=1304400
X182 8498 1 9646 3 505 NAND2X1 $T=1929840 1148560 1 0 $X=1929838 $Y=1143120
X183 9347 1 493 3 9702 NAND2X1 $T=1929840 1269520 0 0 $X=1929838 $Y=1269118
X184 499 1 500 3 9632 NAND2X1 $T=1932480 1350160 0 0 $X=1932478 $Y=1349758
X185 8417 1 9723 3 9738 NAND2X1 $T=1936440 1178800 1 0 $X=1936438 $Y=1173360
X186 435 1 9596 3 9712 NAND2X1 $T=1937760 1279600 0 0 $X=1937758 $Y=1279198
X187 435 1 9667 3 9740 NAND2X1 $T=1940400 1259440 0 0 $X=1940398 $Y=1259038
X188 8575 1 9796 3 9728 NAND2X1 $T=1953600 1209040 1 0 $X=1953598 $Y=1203600
X189 10316 1 10297 3 10330 NAND2X1 $T=2039400 1209040 1 0 $X=2039398 $Y=1203600
X190 10496 1 10432 3 10396 NAND2X1 $T=2051940 1148560 1 180 $X=2049960 $Y=1148158
X191 10572 1 10580 3 10607 NAND2X1 $T=2075700 1330000 0 180 $X=2073720 $Y=1324560
X192 10623 1 10633 3 571 NAND2X1 $T=2085600 1410640 0 0 $X=2085598 $Y=1410238
X193 10702 1 10823 3 10820 NAND2X1 $T=2113980 1380400 1 0 $X=2113978 $Y=1374960
X194 10840 1 10821 3 10868 NAND2X1 $T=2121900 1390480 1 0 $X=2121898 $Y=1385040
X195 10866 1 10865 3 10840 NAND2X1 $T=2123220 1350160 0 0 $X=2123218 $Y=1349758
X196 10883 1 10890 3 10891 NAND2X1 $T=2125860 1420720 1 0 $X=2125858 $Y=1415280
X197 10893 1 10889 3 10883 NAND2X1 $T=2127840 1410640 1 180 $X=2125860 $Y=1410238
X198 10890 1 10863 3 10922 NAND2X1 $T=2131140 1420720 1 0 $X=2131138 $Y=1415280
X199 592 1 11071 3 11094 NAND2X1 $T=2154900 1420720 0 0 $X=2154898 $Y=1420318
X200 11125 1 11259 3 11253 NAND2X1 $T=2189880 1390480 0 0 $X=2189878 $Y=1390078
X201 11182 1 11357 3 11420 NAND2X1 $T=2201760 1330000 1 0 $X=2201758 $Y=1324560
X202 11285 1 11412 3 11445 NAND2X1 $T=2211000 1350160 1 0 $X=2210998 $Y=1344720
X203 11445 1 11454 3 11455 NAND2X1 $T=2219580 1380400 1 180 $X=2217600 $Y=1379998
X204 11356 1 11512 3 11526 NAND2X1 $T=2231460 1309840 0 180 $X=2229480 $Y=1304400
X205 11387 1 11553 3 11555 NAND2X1 $T=2233440 1289680 0 0 $X=2233438 $Y=1289278
X206 11588 1 611 3 11554 NAND2X1 $T=2240700 1390480 1 180 $X=2238720 $Y=1390078
X207 615 1 11738 3 11579 NAND2X1 $T=2266440 1400560 1 180 $X=2264460 $Y=1400158
X208 11905 1 12072 3 12186 NAND2X1 $T=2309340 1148560 0 0 $X=2309338 $Y=1148158
X209 11791 1 11811 3 12126 NAND2X1 $T=2313960 1299760 1 0 $X=2313958 $Y=1294320
X210 11827 1 12165 3 12185 NAND2X1 $T=2324520 1249360 0 0 $X=2324518 $Y=1248958
X211 12132 1 619 3 12041 NAND2X1 $T=2327160 1390480 1 0 $X=2327158 $Y=1385040
X212 11805 1 12159 3 12213 NAND2X1 $T=2329140 1279600 1 0 $X=2329138 $Y=1274160
X213 11826 1 11926 3 12279 NAND2X1 $T=2341680 1209040 1 0 $X=2341678 $Y=1203600
X214 12212 1 11908 3 12325 NAND2X1 $T=2343000 1168720 1 0 $X=2342998 $Y=1163280
X215 12216 1 12288 3 12287 NAND2X1 $T=2344320 1350160 0 0 $X=2344318 $Y=1349758
X216 12275 1 11964 3 12288 NAND2X1 $T=2344320 1360240 0 0 $X=2344318 $Y=1359838
X217 11963 1 11962 3 12286 NAND2X1 $T=2346300 1239280 0 180 $X=2344320 $Y=1233840
X218 12220 1 12131 3 12456 NAND2X1 $T=2349600 1188880 0 0 $X=2349598 $Y=1188478
X219 12213 1 12271 3 12401 NAND2X1 $T=2356860 1279600 0 0 $X=2356858 $Y=1279198
X220 12435 1 12427 3 12326 NAND2X1 $T=2363460 1400560 1 180 $X=2361480 $Y=1400158
X221 12247 1 12398 3 12535 NAND2X1 $T=2369400 1269520 1 0 $X=2369398 $Y=1264080
X222 12271 1 12398 3 12505 NAND2X1 $T=2369400 1279600 0 0 $X=2369398 $Y=1279198
X223 12467 1 12492 3 12522 NAND2X1 $T=2371380 1219120 0 0 $X=2371378 $Y=1218718
X224 12502 1 633 3 12426 NAND2X1 $T=2375340 1350160 1 180 $X=2373360 $Y=1349758
X225 12372 1 12495 3 12466 NAND2X1 $T=2374680 1198960 1 0 $X=2374678 $Y=1193520
X226 12328 1 12503 3 12504 NAND2X1 $T=2376660 1420720 0 0 $X=2376658 $Y=1420318
X227 12456 1 12495 3 12571 NAND2X1 $T=2385900 1198960 0 0 $X=2385898 $Y=1198558
X228 12496 1 12598 3 12560 NAND2X1 $T=2389860 1239280 1 0 $X=2389858 $Y=1233840
X229 12495 1 12622 3 12534 NAND2X1 $T=2393820 1198960 0 0 $X=2393818 $Y=1198558
X230 12492 1 12715 3 12716 NAND2X1 $T=2402400 1229200 0 180 $X=2400420 $Y=1223760
X231 12715 1 12807 3 12774 NAND2X1 $T=2416260 1229200 1 0 $X=2416258 $Y=1223760
X232 12569 1 12770 3 12595 NAND2X1 $T=2421540 1390480 0 0 $X=2421538 $Y=1390078
X233 12628 1 12808 3 12725 NAND2X1 $T=2422860 1370320 0 0 $X=2422858 $Y=1369918
X234 12818 1 12835 3 12935 NAND2X1 $T=2430780 1158640 0 0 $X=2430778 $Y=1158238
X235 12650 1 12888 3 12819 NAND2X1 $T=2442660 1360240 1 0 $X=2442658 $Y=1354800
X236 13116 1 12999 3 12937 NAND2X1 $T=2459820 1319920 1 0 $X=2459818 $Y=1314480
X237 13089 1 13117 3 13124 NAND2X1 $T=2460480 1410640 1 0 $X=2460478 $Y=1405200
X238 13129 1 646 3 13116 NAND2X1 $T=2467740 1330000 1 0 $X=2467738 $Y=1324560
X239 13189 1 13124 3 13180 NAND2X1 $T=2473020 1390480 0 180 $X=2471040 $Y=1385040
X240 12939 1 13218 3 13216 NAND2X1 $T=2476980 1350160 0 0 $X=2476978 $Y=1349758
X241 13305 1 651 3 13272 NAND2X1 $T=2487540 1158640 0 180 $X=2485560 $Y=1153200
X242 654 1 13088 3 13417 NAND2X1 $T=2494800 1420720 0 0 $X=2494798 $Y=1420318
X243 12844 1 13461 3 13500 NAND2X1 $T=2510640 1330000 1 0 $X=2510638 $Y=1324560
X244 13501 1 13207 3 13515 NAND2X1 $T=2512620 1350160 1 0 $X=2512618 $Y=1344720
X245 13317 1 13589 3 13560 NAND2X1 $T=2520540 1198960 0 0 $X=2520538 $Y=1198558
X246 669 1 667 3 13651 NAND2X1 $T=2530440 1420720 1 180 $X=2528460 $Y=1420318
X247 13093 1 13655 3 13610 NAND2X1 $T=2529120 1309840 0 0 $X=2529118 $Y=1309438
X248 13816 1 13684 3 13898 NAND2X1 $T=2548920 1400560 1 180 $X=2546940 $Y=1400158
X249 12722 1 13834 3 13876 NAND2X1 $T=2550900 1259440 0 180 $X=2548920 $Y=1254000
X250 13814 1 13605 3 13835 NAND2X1 $T=2550900 1299760 0 180 $X=2548920 $Y=1294320
X251 671 1 673 3 674 NAND2X1 $T=2549580 1138480 0 0 $X=2549578 $Y=1138078
X252 670 1 672 3 13870 NAND2X1 $T=2549580 1410640 0 0 $X=2549578 $Y=1410238
X253 13876 1 13899 3 13823 NAND2X1 $T=2557500 1259440 0 0 $X=2557498 $Y=1259038
X254 680 1 13900 3 13968 NAND2X1 $T=2559480 1380400 1 180 $X=2557500 $Y=1379998
X255 12870 1 13882 3 13813 NAND2X1 $T=2560800 1309840 1 0 $X=2560798 $Y=1304400
X256 13985 1 13902 3 13937 NAND2X1 $T=2567400 1158640 1 180 $X=2565420 $Y=1158238
X257 13980 1 681 3 13874 NAND2X1 $T=2571360 1188880 1 0 $X=2571358 $Y=1183440
X258 689 1 683 3 14018 NAND2X1 $T=2575320 1430800 0 180 $X=2573340 $Y=1425360
X259 684 1 14020 3 13927 NAND2X1 $T=2575980 1239280 0 0 $X=2575978 $Y=1238878
X260 14035 1 14012 3 14042 NAND2X1 $T=2578620 1279600 0 0 $X=2578618 $Y=1279198
X261 14033 1 14074 3 14072 NAND2X1 $T=2583900 1269520 0 0 $X=2583898 $Y=1269118
X262 690 1 14115 3 14059 NAND2X1 $T=2590500 1168720 1 0 $X=2590498 $Y=1163280
X263 14111 1 13698 3 14074 NAND2X1 $T=2591820 1279600 0 0 $X=2591818 $Y=1279198
X264 14110 1 691 3 14225 NAND2X1 $T=2594460 1370320 1 0 $X=2594458 $Y=1364880
X265 694 1 14227 3 14082 NAND2X1 $T=2601720 1158640 0 0 $X=2601718 $Y=1158238
X266 14139 1 696 3 14257 NAND2X1 $T=2609640 1410640 0 0 $X=2609638 $Y=1410238
X267 12493 1 14279 3 14229 NAND2X1 $T=2612280 1239280 0 0 $X=2612278 $Y=1238878
X268 2140 3 1 2671 2689 NOR2X4 $T=848760 1209040 1 180 $X=844140 $Y=1208638
X269 56 3 1 2875 2870 NOR2X4 $T=875160 1259440 1 180 $X=870540 $Y=1259038
X270 60 3 1 2939 2942 NOR2X4 $T=888360 1340080 0 180 $X=883740 $Y=1334640
X271 116 3 1 2951 2955 NOR2X4 $T=891000 1370320 1 180 $X=886380 $Y=1369918
X272 54 3 1 2949 2956 NOR2X4 $T=891000 1400560 1 180 $X=886380 $Y=1400158
X273 53 3 1 2947 2841 NOR2X4 $T=892320 1289680 1 180 $X=887700 $Y=1289278
X274 59 3 1 3064 3087 NOR2X4 $T=909480 1330000 1 180 $X=904860 $Y=1329598
X275 307 3 1 3379 6339 NOR2X4 $T=1419660 1400560 1 180 $X=1415040 $Y=1400158
X276 2944 3 1 7176 7178 NOR2X4 $T=1547700 1178800 0 180 $X=1543080 $Y=1173360
X277 7391 3 1 2820 7519 NOR2X4 $T=1576740 1158640 1 0 $X=1576738 $Y=1153200
X278 7258 3 1 7597 7598 NOR2X4 $T=1605120 1249360 0 180 $X=1600500 $Y=1243920
X279 7653 3 1 6950 7626 NOR2X4 $T=1610400 1269520 0 180 $X=1605780 $Y=1264080
X280 7982 3 1 7836 7932 NOR2X4 $T=1657260 1168720 1 180 $X=1652640 $Y=1168318
X281 366 3 1 7600 7952 NOR2X4 $T=1662540 1188880 1 180 $X=1657920 $Y=1188478
X282 9002 3 1 8942 9012 NOR2X4 $T=1829520 1370320 1 180 $X=1824900 $Y=1369918
X283 456 3 1 455 9002 NOR2X4 $T=1827540 1390480 1 0 $X=1827538 $Y=1385040
X284 526 3 1 527 9986 NOR2X4 $T=1980000 1370320 1 0 $X=1979998 $Y=1364880
X285 9684 3 1 9985 10003 NOR2X4 $T=1982640 1319920 0 0 $X=1982638 $Y=1319518
X286 529 3 1 530 10036 NOR2X4 $T=1997820 1259440 1 0 $X=1997818 $Y=1254000
X287 537 3 1 536 10236 NOR2X4 $T=2018940 1279600 1 0 $X=2018938 $Y=1274160
X288 540 3 1 539 10264 NOR2X4 $T=2031480 1299760 1 0 $X=2031478 $Y=1294320
X289 616 3 1 11875 11847 NOR2X4 $T=2280300 1410640 1 0 $X=2280298 $Y=1405200
X290 617 3 1 12043 11875 NOR2X4 $T=2304060 1410640 0 0 $X=2304058 $Y=1410238
X291 12502 3 1 633 12399 NOR2X4 $T=2379960 1350160 0 0 $X=2379958 $Y=1349758
X292 13188 3 1 650 13155 NOR2X4 $T=2472360 1289680 1 0 $X=2472358 $Y=1284240
X293 13561 3 1 664 13318 NOR2X4 $T=2518560 1259440 0 0 $X=2518558 $Y=1259038
X294 13701 3 1 668 13609 NOR2X4 $T=2539680 1239280 0 0 $X=2539678 $Y=1238878
X295 13929 3 1 677 13287 NOR2X4 $T=2554200 1209040 0 180 $X=2549580 $Y=1203600
X296 13881 3 1 678 13645 NOR2X4 $T=2560140 1229200 1 0 $X=2560138 $Y=1223760
X297 13980 3 1 681 13785 NOR2X4 $T=2574000 1198960 0 180 $X=2569380 $Y=1193520
X298 77 1 1787 1693 3 NAND2BX1 $T=712140 1430800 0 180 $X=709500 $Y=1425360
X299 1996 1 1989 1775 3 NAND2BX1 $T=741840 1420720 0 180 $X=739200 $Y=1415280
X300 2942 1 2984 2979 3 NAND2BX1 $T=894300 1340080 0 180 $X=891660 $Y=1334640
X301 2955 1 3015 3111 3 NAND2BX1 $T=902220 1370320 0 0 $X=902218 $Y=1369918
X302 3087 1 3022 3172 3 NAND2BX1 $T=920040 1340080 0 0 $X=920038 $Y=1339678
X303 3119 1 3134 3239 3 NAND2BX1 $T=923340 1410640 1 0 $X=923338 $Y=1405200
X304 3270 1 125 3214 3 NAND2BX1 $T=940500 1178800 1 180 $X=937860 $Y=1178398
X305 3404 1 3414 3285 3 NAND2BX1 $T=969540 1239280 1 180 $X=966900 $Y=1238878
X306 3495 1 3481 3466 3 NAND2BX1 $T=977460 1380400 1 180 $X=974820 $Y=1379998
X307 142 1 143 3562 3 NAND2BX1 $T=982740 1148560 1 0 $X=982738 $Y=1143120
X308 150 1 3562 3585 3 NAND2BX1 $T=993300 1148560 0 180 $X=990660 $Y=1143120
X309 3704 1 3699 3586 3 NAND2BX1 $T=1006500 1330000 0 180 $X=1003860 $Y=1324560
X310 3707 1 3698 3703 3 NAND2BX1 $T=1015080 1249360 0 180 $X=1012440 $Y=1243920
X311 3803 1 3804 3815 3 NAND2BX1 $T=1029600 1269520 0 180 $X=1026960 $Y=1264080
X312 3793 1 3866 3702 3 NAND2BX1 $T=1034880 1239280 0 180 $X=1032240 $Y=1233840
X313 4120 1 4090 4053 3 NAND2BX1 $T=1063920 1400560 1 180 $X=1061280 $Y=1400158
X314 4990 1 4958 237 3 NAND2BX1 $T=1207800 1269520 0 180 $X=1205160 $Y=1264080
X315 5276 1 257 5356 3 NAND2BX1 $T=1246740 1239280 1 0 $X=1246738 $Y=1233840
X316 257 1 5276 5375 3 NAND2BX1 $T=1254660 1239280 1 0 $X=1254658 $Y=1233840
X317 6280 1 6279 6310 3 NAND2BX1 $T=1407780 1289680 1 0 $X=1407778 $Y=1284240
X318 6282 1 6281 6426 3 NAND2BX1 $T=1432200 1249360 1 0 $X=1432198 $Y=1243920
X319 6485 1 6630 6724 3 NAND2BX1 $T=1461240 1370320 1 0 $X=1461238 $Y=1364880
X320 6635 1 6575 6762 3 NAND2BX1 $T=1463880 1229200 1 0 $X=1463878 $Y=1223760
X321 6598 1 6660 6661 3 NAND2BX1 $T=1466520 1259440 1 0 $X=1466518 $Y=1254000
X322 6699 1 6732 6795 3 NAND2BX1 $T=1479720 1269520 0 0 $X=1479718 $Y=1269118
X323 6664 1 6735 6837 3 NAND2BX1 $T=1487640 1209040 0 0 $X=1487638 $Y=1208638
X324 7287 1 7378 7387 3 NAND2BX1 $T=1571460 1198960 0 0 $X=1571458 $Y=1198558
X325 7626 1 7650 7698 3 NAND2BX1 $T=1616340 1269520 1 0 $X=1616338 $Y=1264080
X326 7932 1 7981 8073 3 NAND2BX1 $T=1671120 1178800 0 0 $X=1671118 $Y=1178398
X327 8270 1 8266 8305 3 NAND2BX1 $T=1711380 1350160 1 0 $X=1711378 $Y=1344720
X328 8590 1 8622 8632 3 NAND2BX1 $T=1763520 1279600 0 0 $X=1763518 $Y=1279198
X329 9002 1 8981 8951 3 NAND2BX1 $T=1824900 1390480 0 180 $X=1822260 $Y=1385040
X330 9121 1 9101 9075 3 NAND2BX1 $T=1843380 1168720 0 180 $X=1840740 $Y=1163280
X331 9208 1 9190 9077 3 NAND2BX1 $T=1859220 1148560 1 180 $X=1856580 $Y=1148158
X332 9684 1 9814 9894 3 NAND2BX1 $T=1963500 1340080 1 180 $X=1960860 $Y=1339678
X333 9920 1 9814 9957 3 NAND2BX1 $T=1974060 1350160 1 0 $X=1974058 $Y=1344720
X334 10394 1 10357 10232 3 NAND2BX1 $T=2040720 1360240 0 180 $X=2038080 $Y=1354800
X335 10784 1 10820 581 3 NAND2BX1 $T=2112660 1410640 0 0 $X=2112658 $Y=1410238
X336 10860 1 10840 10767 3 NAND2BX1 $T=2120580 1390480 1 180 $X=2117940 $Y=1390078
X337 598 1 11128 11232 3 NAND2BX1 $T=2170080 1430800 1 0 $X=2170078 $Y=1425360
X338 11251 1 11253 603 3 NAND2BX1 $T=2188560 1400560 0 0 $X=2188558 $Y=1400158
X339 11585 1 11555 11705 3 NAND2BX1 $T=2247300 1319920 1 0 $X=2247298 $Y=1314480
X340 12221 1 12216 12074 3 NAND2BX1 $T=2333100 1360240 0 180 $X=2330460 $Y=1354800
X341 12270 1 12276 12324 3 NAND2BX1 $T=2341680 1148560 1 0 $X=2341678 $Y=1143120
X342 12397 1 12326 12245 3 NAND2BX1 $T=2350920 1400560 1 180 $X=2348280 $Y=1400158
X343 12130 1 12186 12568 3 NAND2BX1 $T=2384580 1158640 1 0 $X=2384578 $Y=1153200
X344 12477 1 12595 12322 3 NAND2BX1 $T=2391180 1390480 1 180 $X=2388540 $Y=1390078
X345 12535 1 12496 12624 3 NAND2BX1 $T=2392500 1239280 0 0 $X=2392498 $Y=1238878
X346 12717 1 12725 12633 3 NAND2BX1 $T=2408340 1370320 1 180 $X=2405700 $Y=1369918
X347 12777 1 12819 12744 3 NAND2BX1 $T=2421540 1360240 0 180 $X=2418900 $Y=1354800
X348 13318 1 13348 13246 3 NAND2BX1 $T=2512620 1259440 1 180 $X=2509980 $Y=1259038
X349 13645 1 13638 13419 3 NAND2BX1 $T=2528460 1229200 0 180 $X=2525820 $Y=1223760
X350 13812 1 13790 13765 3 NAND2BX1 $T=2548260 1148560 1 180 $X=2545620 $Y=1148158
X351 13971 1 13968 13986 3 NAND2BX1 $T=2570040 1360240 0 0 $X=2570038 $Y=1359838
X352 13898 1 683 14041 3 NAND2BX1 $T=2580600 1410640 1 0 $X=2580598 $Y=1405200
X353 14071 1 14059 14046 3 NAND2BX1 $T=2583240 1178800 1 180 $X=2580600 $Y=1178398
X354 13975 1 14088 14060 3 NAND2BX1 $T=2585880 1259440 0 0 $X=2585878 $Y=1259038
X355 1840 55 1 1886 3 1889 OAI21X1 $T=723360 1249360 1 0 $X=723358 $Y=1243920
X356 1956 1916 1 1958 3 1954 OAI21X1 $T=733920 1360240 1 0 $X=733918 $Y=1354800
X357 3803 3801 1 3804 3 3749 OAI21X1 $T=1021680 1259440 0 0 $X=1021678 $Y=1259038
X358 3699 3812 1 3836 3 3750 OAI21X1 $T=1024320 1319920 0 0 $X=1024318 $Y=1319518
X359 6281 6307 1 6306 3 6308 OAI21X1 $T=1412400 1239280 0 180 $X=1409100 $Y=1233840
X360 6255 6280 1 6279 3 6457 OAI21X1 $T=1414380 1289680 1 0 $X=1414378 $Y=1284240
X361 8892 8882 1 8862 3 8792 OAI21X1 $T=1805100 1168720 0 180 $X=1801800 $Y=1163280
X362 8887 8883 1 8892 3 8940 OAI21X1 $T=1813020 1188880 1 0 $X=1813018 $Y=1183440
X363 9732 9703 1 9668 3 9627 OAI21X1 $T=1932480 1330000 1 180 $X=1929180 $Y=1329598
X364 10922 579 1 10945 3 11092 OAI21X1 $T=2136420 1420720 1 0 $X=2136418 $Y=1415280
X365 11251 11179 1 11253 3 11279 OAI21X1 $T=2186580 1410640 0 0 $X=2186578 $Y=1410238
X366 11445 11417 1 11420 3 11444 OAI21X1 $T=2217600 1340080 0 180 $X=2214300 $Y=1334640
X367 11546 11578 1 11526 3 11582 OAI21X1 $T=2241360 1360240 0 180 $X=2238060 $Y=1354800
X368 12213 12246 1 12185 3 12374 OAI21X1 $T=2346300 1269520 1 0 $X=2346298 $Y=1264080
X369 12130 634 1 12186 3 12649 OAI21X1 $T=2382600 1148560 1 0 $X=2382598 $Y=1143120
X370 12624 12192 1 12599 3 12602 OAI21X1 $T=2393160 1249360 1 180 $X=2389860 $Y=1248958
X371 12716 12192 1 12721 3 12802 OAI21X1 $T=2401080 1239280 0 0 $X=2401078 $Y=1238878
X372 13835 13508 1 13808 3 13807 OAI21X1 $T=2550900 1279600 1 180 $X=2547600 $Y=1279198
X373 13424 13785 1 13874 3 13691 OAI21X1 $T=2550240 1188880 0 0 $X=2550238 $Y=1188478
X374 13808 14060 1 14224 3 14118 OAI21X1 $T=2597760 1269520 0 0 $X=2597758 $Y=1269118
X375 1545 1 67 1572 3 1569 OAI21XL $T=677820 1289680 1 0 $X=677818 $Y=1284240
X376 1603 1 1574 1576 3 1577 OAI21XL $T=683100 1219120 0 180 $X=680460 $Y=1213680
X377 1609 1 55 1629 3 1571 OAI21XL $T=684420 1249360 0 180 $X=681780 $Y=1243920
X378 1605 1 1657 1603 3 1656 OAI21XL $T=693660 1239280 1 180 $X=691020 $Y=1238878
X379 1754 1 76 1778 3 1776 OAI21XL $T=705540 1350160 0 0 $X=705538 $Y=1349758
X380 1849 1 76 1821 3 1774 OAI21XL $T=718080 1410640 1 180 $X=715440 $Y=1410238
X381 1898 1 76 1916 3 1919 OAI21XL $T=726660 1400560 0 0 $X=726658 $Y=1400158
X382 2138 1 1986 2135 3 2107 OAI21XL $T=752400 1168720 1 180 $X=749760 $Y=1168318
X383 1841 1 2142 2145 3 2111 OAI21XL $T=759000 1340080 1 180 $X=756360 $Y=1339678
X384 1917 1 1996 1989 3 2018 OAI21XL $T=757680 1420720 1 0 $X=757678 $Y=1415280
X385 2170 1 1986 2278 3 2115 OAI21XL $T=762960 1219120 0 180 $X=760320 $Y=1213680
X386 2172 1 1986 2181 3 2137 OAI21XL $T=763620 1279600 1 0 $X=763618 $Y=1274160
X387 1980 1 2113 2167 3 1752 OAI21XL $T=766260 1370320 1 180 $X=763620 $Y=1369918
X388 2214 1 2207 2202 3 2139 OAI21XL $T=768240 1168720 0 180 $X=765600 $Y=1163280
X389 2211 1 1986 2243 3 2180 OAI21XL $T=768900 1249360 0 180 $X=766260 $Y=1243920
X390 2215 1 1986 2235 3 2157 OAI21XL $T=769560 1299760 1 0 $X=769558 $Y=1294320
X391 2251 1 1986 2207 3 2299 OAI21XL $T=774840 1168720 0 0 $X=774838 $Y=1168318
X392 2281 1 2235 2285 3 2276 OAI21XL $T=778800 1279600 1 0 $X=778798 $Y=1274160
X393 2235 1 2237 2317 3 2270 OAI21XL $T=782760 1269520 1 0 $X=782758 $Y=1264080
X394 2368 1 1986 2349 3 2350 OAI21XL $T=792000 1188880 0 0 $X=791998 $Y=1188478
X395 2285 1 2321 2346 3 2386 OAI21XL $T=794640 1279600 1 0 $X=794638 $Y=1274160
X396 3273 1 3404 3414 3 3354 OAI21XL $T=961620 1239280 0 0 $X=961618 $Y=1238878
X397 3478 1 3475 3465 3 3412 OAI21XL $T=974820 1299760 0 180 $X=972180 $Y=1294320
X398 3434 1 3437 3478 3 3252 OAI21XL $T=976140 1309840 0 180 $X=973500 $Y=1304400
X399 3704 1 3672 3699 3 3673 OAI21XL $T=1006500 1340080 0 180 $X=1003860 $Y=1334640
X400 3615 1 3694 3711 3 150 OAI21XL $T=1007160 1168720 0 0 $X=1007158 $Y=1168318
X401 3698 1 3793 3866 3 3744 OAI21XL $T=1032240 1229200 0 0 $X=1032238 $Y=1228798
X402 208 1 4666 4669 3 220 OAI21XL $T=1164240 1188880 0 180 $X=1161600 $Y=1183440
X403 219 1 192 4617 3 4722 OAI21XL $T=1164240 1370320 1 0 $X=1164238 $Y=1364880
X404 4666 1 189 4669 3 5063 OAI21XL $T=1169520 1188880 0 0 $X=1169518 $Y=1188478
X405 4724 1 4722 4670 3 4851 OAI21XL $T=1172160 1370320 1 0 $X=1172158 $Y=1364880
X406 218 1 230 4785 3 227 OAI21XL $T=1186020 1168720 1 180 $X=1183380 $Y=1168318
X407 222 1 4814 4720 3 4881 OAI21XL $T=1188000 1380400 0 0 $X=1187998 $Y=1379998
X408 232 1 192 204 3 4785 OAI21XL $T=1195920 1168720 1 180 $X=1193280 $Y=1168318
X409 210 1 232 221 3 4885 OAI21XL $T=1201200 1249360 1 180 $X=1198560 $Y=1248958
X410 230 1 191 4885 3 4891 OAI21XL $T=1202520 1239280 0 180 $X=1199880 $Y=1233840
X411 4953 1 4947 4952 3 4955 OAI21XL $T=1203840 1209040 1 0 $X=1203838 $Y=1203600
X412 210 1 230 228 3 4958 OAI21XL $T=1203840 1259440 0 0 $X=1203838 $Y=1259038
X413 5022 1 192 5019 3 4952 OAI21XL $T=1206480 1229200 1 180 $X=1203840 $Y=1228798
X414 4778 1 192 4849 3 243 OAI21XL $T=1205160 1138480 0 0 $X=1205158 $Y=1138078
X415 5063 1 4954 199 3 5102 OAI21XL $T=1219680 1188880 0 0 $X=1219678 $Y=1188478
X416 4954 1 5022 5019 3 5354 OAI21XL $T=1228260 1229200 0 0 $X=1228258 $Y=1228798
X417 246 1 189 5103 3 5213 OAI21XL $T=1228260 1410640 1 0 $X=1228258 $Y=1405200
X418 5072 1 5109 5135 3 5192 OAI21XL $T=1234860 1289680 1 0 $X=1234858 $Y=1284240
X419 5198 1 5213 5143 3 5222 OAI21XL $T=1237500 1400560 0 0 $X=1237498 $Y=1400158
X420 5233 1 253 5237 3 5221 OAI21XL $T=1241460 1259440 1 180 $X=1238820 $Y=1259038
X421 4990 1 5234 5227 3 5237 OAI21XL $T=1240140 1269520 1 0 $X=1240138 $Y=1264080
X422 247 1 187 5226 3 5304 OAI21XL $T=1242780 1198960 0 0 $X=1242778 $Y=1198558
X423 5262 1 5264 253 3 5345 OAI21XL $T=1243440 1168720 1 0 $X=1243438 $Y=1163280
X424 4954 1 5185 5266 3 5276 OAI21XL $T=1244100 1239280 0 0 $X=1244098 $Y=1238878
X425 5226 1 5303 204 3 5346 OAI21XL $T=1253340 1198960 1 180 $X=1250700 $Y=1198558
X426 5520 1 5542 5220 3 5584 OAI21XL $T=1287000 1178800 0 0 $X=1286998 $Y=1178398
X427 5553 1 5488 5487 3 5675 OAI21XL $T=1310760 1148560 0 0 $X=1310758 $Y=1148158
X428 5948 1 128 5944 3 5972 OAI21XL $T=1359600 1420720 1 0 $X=1359598 $Y=1415280
X429 6002 1 134 5998 3 5999 OAI21XL $T=1369500 1400560 1 180 $X=1366860 $Y=1400158
X430 5999 1 6029 6030 3 6038 OAI21XL $T=1369500 1410640 1 0 $X=1369498 $Y=1405200
X431 6002 1 200 6001 3 6250 OAI21XL $T=1378740 1370320 0 0 $X=1378738 $Y=1369918
X432 6250 1 6193 6040 3 6256 OAI21XL $T=1399860 1370320 0 0 $X=1399858 $Y=1369918
X433 5948 1 197 6190 3 6365 OAI21XL $T=1415040 1390480 1 0 $X=1415038 $Y=1385040
X434 7138 1 6998 335 3 7259 OAI21XL $T=1550340 1289680 1 0 $X=1550338 $Y=1284240
X435 7282 1 6998 7283 3 7263 OAI21XL $T=1558260 1239280 1 180 $X=1555620 $Y=1238878
X436 7321 1 7266 7278 3 7390 OAI21XL $T=1562220 1350160 1 0 $X=1562218 $Y=1344720
X437 7261 1 7266 7214 3 7353 OAI21XL $T=1564200 1370320 1 0 $X=1564198 $Y=1364880
X438 7626 1 7677 7650 3 7719 OAI21XL $T=1618320 1259440 0 0 $X=1618318 $Y=1259038
X439 376 1 368 375 3 8120 OAI21XL $T=1691580 1390480 1 180 $X=1688940 $Y=1390078
X440 8150 1 8270 8266 3 8264 OAI21XL $T=1706100 1340080 1 0 $X=1706098 $Y=1334640
X441 8860 1 8859 8861 3 8865 OAI21XL $T=1806420 1370320 0 180 $X=1803780 $Y=1364880
X442 8942 1 8859 8945 3 8948 OAI21XL $T=1815660 1370320 0 0 $X=1815658 $Y=1369918
X443 9121 1 9074 9101 3 9073 OAI21XL $T=1847340 1158640 0 180 $X=1844700 $Y=1153200
X444 9187 1 479 9204 3 482 OAI21XL $T=1877700 1430800 1 0 $X=1877698 $Y=1425360
X445 487 1 9441 488 3 490 OAI21XL $T=1896840 1430800 1 0 $X=1896838 $Y=1425360
X446 10323 1 10318 10330 3 10329 OAI21XL $T=2034120 1198960 1 0 $X=2034118 $Y=1193520
X447 534 1 10394 10357 3 10392 OAI21XL $T=2048640 1360240 0 180 $X=2046000 $Y=1354800
X448 10621 1 10617 10607 3 10609 OAI21XL $T=2083620 1330000 0 180 $X=2080980 $Y=1324560
X449 11232 1 601 11179 3 602 OAI21XL $T=2185920 1420720 0 0 $X=2185918 $Y=1420318
X450 11526 1 11585 11555 3 11599 OAI21XL $T=2239380 1309840 0 0 $X=2239378 $Y=1309438
X451 12186 1 12270 12276 3 628 OAI21XL $T=2350260 1148560 1 0 $X=2350258 $Y=1143120
X452 12292 1 12466 12460 3 12433 OAI21XL $T=2370060 1198960 0 180 $X=2367420 $Y=1193520
X453 12535 1 12192 12436 3 12559 OAI21XL $T=2386560 1269520 0 180 $X=2383920 $Y=1264080
X454 12774 1 12192 12778 3 12817 OAI21XL $T=2410980 1239280 1 0 $X=2410978 $Y=1233840
X455 12903 1 634 12895 3 13128 OAI21XL $T=2434080 1158640 1 0 $X=2434078 $Y=1153200
X456 12909 1 634 12904 3 12956 OAI21XL $T=2439360 1148560 1 0 $X=2439358 $Y=1143120
X457 642 1 643 644 3 12978 OAI21XL $T=2443320 1420720 0 0 $X=2443318 $Y=1420318
X458 648 1 644 649 3 13179 OAI21XL $T=2472360 1430800 1 0 $X=2472358 $Y=1425360
X459 660 1 13308 661 3 13516 OAI21XL $T=2504700 1410640 0 0 $X=2504698 $Y=1410238
X460 13417 1 643 13428 3 13433 OAI21XL $T=2505360 1420720 0 0 $X=2505358 $Y=1420318
X461 13562 1 643 13520 3 13525 OAI21XL $T=2517900 1410640 0 180 $X=2515260 $Y=1405200
X462 13743 1 13219 13651 3 13815 OAI21XL $T=2540340 1400560 1 0 $X=2540338 $Y=1395120
X463 674 1 13812 13790 3 13885 OAI21XL $T=2553540 1148560 0 0 $X=2553538 $Y=1148158
X464 13913 1 13219 13912 3 13869 OAI21XL $T=2561460 1370320 0 180 $X=2558820 $Y=1364880
X465 13941 1 13937 13906 3 13286 OAI21XL $T=2562120 1158640 1 180 $X=2559480 $Y=1158238
X466 13898 1 13219 13877 3 13951 OAI21XL $T=2560140 1410640 1 0 $X=2560138 $Y=1405200
X467 13941 1 13949 13945 3 13763 OAI21XL $T=2567400 1138480 1 180 $X=2564760 $Y=1138078
X468 13971 1 13972 13968 3 13931 OAI21XL $T=2570040 1380400 0 180 $X=2567400 $Y=1374960
X469 14018 1 13877 685 3 14010 OAI21XL $T=2576640 1420720 0 180 $X=2574000 $Y=1415280
X470 14076 1 13941 14050 3 686 OAI21XL $T=2580600 1148560 0 180 $X=2577960 $Y=1143120
X471 14011 1 13876 13927 3 14021 OAI21XL $T=2583240 1259440 0 180 $X=2580600 $Y=1254000
X472 13987 1 13219 13972 3 13981 OAI21XL $T=2583240 1370320 0 180 $X=2580600 $Y=1364880
X473 14059 1 14064 14082 3 13950 OAI21XL $T=2584560 1158640 1 0 $X=2584558 $Y=1153200
X474 14228 1 14226 14225 3 14161 OAI21XL $T=2603040 1370320 0 180 $X=2600400 $Y=1364880
X475 13927 1 14073 14229 3 14283 OAI21XL $T=2601720 1249360 1 0 $X=2601718 $Y=1243920
X476 14312 1 13219 14334 3 14127 OAI21XL $T=2618880 1400560 0 0 $X=2618878 $Y=1400158
X477 14338 1 13219 14277 3 14335 OAI21XL $T=2625480 1370320 1 0 $X=2625478 $Y=1364880
X478 1568 1596 71 1 3 XOR2X4 $T=677820 1188880 0 0 $X=677818 $Y=1188478
X479 1914 1925 2171 1 3 XOR2X4 $T=727320 1198960 0 0 $X=727318 $Y=1198558
X480 1981 1564 2140 1 3 XOR2X4 $T=739200 1249360 0 0 $X=739198 $Y=1248958
X481 2986 2978 3093 1 3 XOR2X4 $T=894960 1309840 1 0 $X=894958 $Y=1304400
X482 3108 2954 3274 1 3 XOR2X4 $T=912120 1269520 0 0 $X=912118 $Y=1269118
X483 3172 3156 3352 1 3 XOR2X4 $T=927300 1340080 0 0 $X=927298 $Y=1339678
X484 123 124 3224 1 3 XOR2X4 $T=927300 1430800 1 0 $X=927298 $Y=1425360
X485 3269 3236 3064 1 3 XOR2X4 $T=945120 1319920 0 180 $X=933900 $Y=1314480
X486 3239 3184 3379 1 3 XOR2X4 $T=937860 1400560 0 0 $X=937858 $Y=1400158
X487 106 5486 268 1 3 XOR2X4 $T=1269840 1319920 0 0 $X=1269838 $Y=1319518
X488 279 5654 283 1 3 XOR2X4 $T=1306800 1249360 1 0 $X=1306798 $Y=1243920
X489 282 284 288 1 3 XOR2X4 $T=1322640 1360240 1 0 $X=1322638 $Y=1354800
X490 108 5586 291 1 3 XOR2X4 $T=1328580 1198960 0 0 $X=1328578 $Y=1198558
X491 6567 6599 6629 1 3 XOR2X4 $T=1450680 1168720 0 0 $X=1450678 $Y=1168318
X492 6820 7001 7177 1 3 XOR2X4 $T=1510740 1319920 0 0 $X=1510738 $Y=1319518
X493 7030 7166 7288 1 3 XOR2X4 $T=1539120 1229200 1 0 $X=1539118 $Y=1223760
X494 7387 7632 7655 1 3 XOR2X4 $T=1604460 1188880 0 0 $X=1604458 $Y=1188478
X495 7675 7624 7836 1 3 XOR2X4 $T=1617000 1168720 0 0 $X=1616998 $Y=1168318
X496 470 9692 525 1 3 XOR2X4 $T=1927860 1380400 0 0 $X=1927858 $Y=1379998
X497 516 10421 559 1 3 XOR2X4 $T=2049300 1390480 0 0 $X=2049298 $Y=1390078
X498 11762 11703 7162 1 3 XOR2X4 $T=2257200 1410640 1 180 $X=2245980 $Y=1410238
X499 11874 11844 7256 1 3 XOR2X4 $T=2282940 1380400 1 180 $X=2271720 $Y=1379998
X500 12629 12600 7502 1 3 XOR2X4 $T=2397780 1319920 1 180 $X=2386560 $Y=1319518
X501 12937 12902 12876 1 3 XOR2X4 $T=2440020 1309840 1 180 $X=2428800 $Y=1309438
X502 13245 13222 7806 1 3 XOR2X4 $T=2486880 1198960 1 180 $X=2475660 $Y=1198558
X503 13273 13269 7982 1 3 XOR2X4 $T=2493480 1178800 1 180 $X=2482260 $Y=1178398
X504 14138 14108 13980 1 3 XOR2X4 $T=2597100 1188880 1 180 $X=2585880 $Y=1188478
X505 1509 1 3 1566 INVX1 $T=674520 1249360 1 0 $X=674518 $Y=1243920
X506 1599 1 3 1612 INVX1 $T=686400 1319920 1 0 $X=686398 $Y=1314480
X507 1658 1 3 1660 INVX1 $T=692340 1370320 0 0 $X=692338 $Y=1369918
X508 1744 1 3 1657 INVX1 $T=702240 1259440 1 180 $X=700920 $Y=1259038
X509 1746 1 3 1669 INVX1 $T=702240 1380400 1 180 $X=700920 $Y=1379998
X510 1898 1 3 1750 INVX1 $T=712800 1370320 1 180 $X=711480 $Y=1369918
X511 1839 1 3 1870 INVX1 $T=716760 1279600 1 0 $X=716758 $Y=1274160
X512 1916 1 3 1807 INVX1 $T=722700 1370320 0 180 $X=721380 $Y=1364880
X513 1915 1 3 1885 INVX1 $T=729300 1259440 1 0 $X=729298 $Y=1254000
X514 2166 1 3 1848 INVX1 $T=746460 1350160 0 180 $X=745140 $Y=1344720
X515 2139 1 3 2135 INVX1 $T=757020 1168720 0 180 $X=755700 $Y=1163280
X516 2215 1 3 2110 INVX1 $T=767580 1289680 0 180 $X=766260 $Y=1284240
X517 2212 1 3 2211 INVX1 $T=775500 1249360 0 180 $X=774180 $Y=1243920
X518 2276 1 3 2181 INVX1 $T=775500 1279600 0 180 $X=774180 $Y=1274160
X519 2281 1 3 2177 INVX1 $T=778140 1279600 1 180 $X=776820 $Y=1279198
X520 2275 1 3 2279 INVX1 $T=779460 1229200 0 0 $X=779458 $Y=1228798
X521 2270 1 3 2243 INVX1 $T=780780 1249360 0 180 $X=779460 $Y=1243920
X522 2302 1 3 2316 INVX1 $T=784740 1188880 1 0 $X=784738 $Y=1183440
X523 2353 1 3 2323 INVX1 $T=791340 1198960 0 180 $X=790020 $Y=1193520
X524 2386 1 3 2317 INVX1 $T=796620 1269520 0 180 $X=795300 $Y=1264080
X525 87 1 3 91 INVX1 $T=796620 1360240 1 180 $X=795300 $Y=1359838
X526 103 1 3 2512 INVX1 $T=818400 1289680 0 0 $X=818398 $Y=1289278
X527 2642 1 3 2761 INVX1 $T=842160 1188880 1 0 $X=842158 $Y=1183440
X528 2689 1 3 2766 INVX1 $T=854040 1209040 1 180 $X=852720 $Y=1208638
X529 2872 1 3 2874 INVX1 $T=871860 1178800 1 0 $X=871858 $Y=1173360
X530 2842 1 3 2977 INVX1 $T=886380 1209040 0 0 $X=886378 $Y=1208638
X531 120 1 3 3059 INVX1 $T=909480 1148560 1 0 $X=909478 $Y=1143120
X532 121 1 3 3020 INVX1 $T=916740 1148560 0 180 $X=915420 $Y=1143120
X533 3134 1 3 3089 INVX1 $T=917400 1390480 0 0 $X=917398 $Y=1390078
X534 3069 1 3 3161 INVX1 $T=918060 1380400 0 0 $X=918058 $Y=1379998
X535 3197 1 3 3160 INVX1 $T=932580 1148560 1 180 $X=931260 $Y=1148158
X536 3214 1 3 3142 INVX1 $T=935220 1178800 0 180 $X=933900 $Y=1173360
X537 3264 1 3 3216 INVX1 $T=942480 1299760 0 180 $X=941160 $Y=1294320
X538 3266 1 3 3270 INVX1 $T=945120 1178800 1 180 $X=943800 $Y=1178398
X539 3435 1 3 3419 INVX1 $T=974160 1350160 1 180 $X=972840 $Y=1349758
X540 3586 1 3 3588 INVX1 $T=991320 1340080 0 0 $X=991318 $Y=1339678
X541 3708 1 3 3672 INVX1 $T=1013100 1340080 1 180 $X=1011780 $Y=1339678
X542 167 1 3 3674 INVX1 $T=1026300 1148560 0 180 $X=1024980 $Y=1143120
X543 3898 1 3 3900 INVX1 $T=1036860 1360240 1 0 $X=1036858 $Y=1354800
X544 3924 1 3 3854 INVX1 $T=1042140 1279600 1 180 $X=1040820 $Y=1279198
X545 3955 1 3 3861 INVX1 $T=1044780 1380400 0 180 $X=1043460 $Y=1374960
X546 4090 1 3 4028 INVX1 $T=1065900 1390480 1 180 $X=1064580 $Y=1390078
X547 4120 1 3 4050 INVX1 $T=1068540 1400560 1 180 $X=1067220 $Y=1400158
X548 175 1 3 4126 INVX1 $T=1074480 1420720 1 180 $X=1073160 $Y=1420318
X549 193 1 3 4269 INVX1 $T=1102200 1269520 1 180 $X=1100880 $Y=1269118
X550 4451 1 3 190 INVX1 $T=1112760 1430800 0 180 $X=1111440 $Y=1425360
X551 183 1 3 4367 INVX1 $T=1112760 1299760 0 0 $X=1112758 $Y=1299358
X552 213 1 3 4615 INVX1 $T=1145760 1370320 1 0 $X=1145758 $Y=1364880
X553 4434 1 3 219 INVX1 $T=1153020 1380400 1 0 $X=1153018 $Y=1374960
X554 221 1 3 4307 INVX1 $T=1170180 1390480 1 180 $X=1168860 $Y=1390078
X555 206 1 3 4725 INVX1 $T=1176120 1380400 1 180 $X=1174800 $Y=1379998
X556 198 1 3 4459 INVX1 $T=1183380 1219120 1 180 $X=1182060 $Y=1218718
X557 223 1 3 222 INVX1 $T=1184700 1400560 1 0 $X=1184698 $Y=1395120
X558 221 1 3 4844 INVX1 $T=1191960 1209040 0 0 $X=1191958 $Y=1208638
X559 4890 1 3 4957 INVX1 $T=1200540 1168720 0 0 $X=1200538 $Y=1168318
X560 4988 1 3 4949 INVX1 $T=1209780 1350160 0 180 $X=1208460 $Y=1344720
X561 4891 1 3 5264 INVX1 $T=1221000 1168720 0 0 $X=1220998 $Y=1168318
X562 5099 1 3 246 INVX1 $T=1222320 1410640 0 180 $X=1221000 $Y=1405200
X563 247 1 3 249 INVX1 $T=1224960 1319920 0 180 $X=1223640 $Y=1314480
X564 4990 1 3 5233 INVX1 $T=1231560 1269520 1 0 $X=1231558 $Y=1264080
X565 188 1 3 4954 INVX1 $T=1233540 1239280 0 0 $X=1233538 $Y=1238878
X566 5192 1 3 5227 INVX1 $T=1236840 1279600 0 0 $X=1236838 $Y=1279198
X567 253 1 3 5234 INVX1 $T=1248720 1269520 0 180 $X=1247400 $Y=1264080
X568 5347 1 3 5305 INVX1 $T=1251360 1400560 0 180 $X=1250040 $Y=1395120
X569 252 1 3 255 INVX1 $T=1251360 1410640 1 180 $X=1250040 $Y=1410238
X570 258 1 3 256 INVX1 $T=1251360 1420720 1 180 $X=1250040 $Y=1420318
X571 5262 1 3 5353 INVX1 $T=1252680 1168720 1 0 $X=1252678 $Y=1163280
X572 5264 1 3 5376 INVX1 $T=1257960 1158640 0 0 $X=1257958 $Y=1158238
X573 4811 1 3 5373 INVX1 $T=1257960 1219120 1 0 $X=1257958 $Y=1213680
X574 5350 1 3 5489 INVX1 $T=1268520 1158640 1 0 $X=1268518 $Y=1153200
X575 5304 1 3 5463 INVX1 $T=1274460 1198960 0 0 $X=1274458 $Y=1198558
X576 5433 1 3 5485 INVX1 $T=1278420 1158640 1 0 $X=1278418 $Y=1153200
X577 5492 1 3 5614 INVX1 $T=1280400 1289680 1 0 $X=1280398 $Y=1284240
X578 5411 1 3 5649 INVX1 $T=1284360 1249360 0 0 $X=1284358 $Y=1248958
X579 5542 1 3 5605 INVX1 $T=1288980 1168720 0 0 $X=1288978 $Y=1168318
X580 5463 1 3 5548 INVX1 $T=1289640 1209040 0 0 $X=1289638 $Y=1208638
X581 5520 1 3 5650 INVX1 $T=1302840 1178800 0 0 $X=1302838 $Y=1178398
X582 5348 1 3 5711 INVX1 $T=1307460 1279600 1 0 $X=1307458 $Y=1274160
X583 179 1 3 289 INVX1 $T=1318680 1410640 0 0 $X=1318678 $Y=1410238
X584 5588 1 3 6005 INVX1 $T=1321980 1219120 1 0 $X=1321978 $Y=1213680
X585 5742 1 3 293 INVX1 $T=1350360 1158640 1 0 $X=1350358 $Y=1153200
X586 5673 1 3 5994 INVX1 $T=1353660 1188880 1 0 $X=1353658 $Y=1183440
X587 5781 1 3 5997 INVX1 $T=1354320 1330000 1 0 $X=1354318 $Y=1324560
X588 5810 1 3 6068 INVX1 $T=1362900 1319920 1 0 $X=1362898 $Y=1314480
X589 5925 1 3 5923 INVX1 $T=1364220 1360240 0 0 $X=1364218 $Y=1359838
X590 6038 1 3 6066 INVX1 $T=1375440 1410640 1 0 $X=1375438 $Y=1405200
X591 6099 1 3 6128 INVX1 $T=1383360 1340080 1 0 $X=1383358 $Y=1334640
X592 303 1 3 6123 INVX1 $T=1396560 1390480 1 180 $X=1395240 $Y=1390078
X593 303 1 3 5849 INVX1 $T=1397880 1410640 0 180 $X=1396560 $Y=1405200
X594 304 1 3 5948 INVX1 $T=1397880 1420720 0 180 $X=1396560 $Y=1415280
X595 6192 1 3 6254 INVX1 $T=1398540 1319920 1 0 $X=1398538 $Y=1314480
X596 6256 1 3 6343 INVX1 $T=1412400 1370320 0 0 $X=1412398 $Y=1369918
X597 6278 1 3 6402 INVX1 $T=1417020 1188880 1 0 $X=1417018 $Y=1183440
X598 6368 1 3 6428 INVX1 $T=1432860 1178800 0 0 $X=1432858 $Y=1178398
X599 6282 1 3 6432 INVX1 $T=1433520 1239280 0 0 $X=1433518 $Y=1238878
X600 6433 1 3 6566 INVX1 $T=1440780 1279600 1 0 $X=1440778 $Y=1274160
X601 6423 1 3 6505 INVX1 $T=1446060 1209040 1 0 $X=1446058 $Y=1203600
X602 6459 1 3 6597 INVX1 $T=1448700 1410640 1 0 $X=1448698 $Y=1405200
X603 314 1 3 6002 INVX1 $T=1452660 1370320 1 180 $X=1451340 $Y=1369918
X604 6004 1 3 6693 INVX1 $T=1453980 1158640 1 0 $X=1453978 $Y=1153200
X605 6593 1 3 6632 INVX1 $T=1455300 1340080 0 0 $X=1455298 $Y=1339678
X606 6434 1 3 6628 INVX1 $T=1456620 1410640 1 0 $X=1456618 $Y=1405200
X607 312 1 3 6704 INVX1 $T=1469820 1400560 1 0 $X=1469818 $Y=1395120
X608 6763 1 3 6847 INVX1 $T=1483020 1330000 1 0 $X=1483018 $Y=1324560
X609 6792 1 3 6790 INVX1 $T=1488960 1168720 1 180 $X=1487640 $Y=1168318
X610 6752 1 3 6836 INVX1 $T=1488300 1158640 1 0 $X=1488298 $Y=1153200
X611 6796 1 3 6868 INVX1 $T=1490280 1299760 0 0 $X=1490278 $Y=1299358
X612 6768 1 3 6769 INVX1 $T=1492920 1229200 0 0 $X=1492918 $Y=1228798
X613 325 1 3 6028 INVX1 $T=1497540 1390480 0 180 $X=1496220 $Y=1385040
X614 6940 1 3 6841 INVX1 $T=1506120 1330000 0 0 $X=1506118 $Y=1329598
X615 6798 1 3 6976 INVX1 $T=1506120 1350160 1 0 $X=1506118 $Y=1344720
X616 329 1 3 6878 INVX1 $T=1506120 1400560 0 0 $X=1506118 $Y=1400158
X617 334 1 3 7036 INVX1 $T=1524600 1289680 0 0 $X=1524598 $Y=1289278
X618 7028 1 3 7088 INVX1 $T=1527240 1229200 1 0 $X=1527238 $Y=1223760
X619 7056 1 3 7065 INVX1 $T=1527240 1400560 0 0 $X=1527238 $Y=1400158
X620 333 1 3 7094 INVX1 $T=1529880 1138480 0 0 $X=1529878 $Y=1138078
X621 7073 1 3 7133 INVX1 $T=1535160 1390480 1 0 $X=1535158 $Y=1385040
X622 7129 1 3 7138 INVX1 $T=1540440 1289680 1 0 $X=1540438 $Y=1284240
X623 7074 1 3 7257 INVX1 $T=1540440 1350160 0 0 $X=1540438 $Y=1349758
X624 7214 1 3 7260 INVX1 $T=1552980 1370320 1 0 $X=1552978 $Y=1364880
X625 337 1 3 7265 INVX1 $T=1557600 1289680 1 180 $X=1556280 $Y=1289278
X626 338 1 3 7289 INVX1 $T=1560240 1259440 0 180 $X=1558920 $Y=1254000
X627 7255 1 3 7381 INVX1 $T=1563540 1178800 1 0 $X=1563538 $Y=1173360
X628 7378 1 3 7386 INVX1 $T=1578060 1188880 1 180 $X=1576740 $Y=1188478
X629 7261 1 3 7292 INVX1 $T=1579380 1370320 0 0 $X=1579378 $Y=1369918
X630 345 1 3 7466 INVX1 $T=1590600 1420720 1 180 $X=1589280 $Y=1420318
X631 7471 1 3 7511 INVX1 $T=1589940 1299760 1 0 $X=1589938 $Y=1294320
X632 344 1 3 7415 INVX1 $T=1593900 1239280 1 180 $X=1592580 $Y=1238878
X633 7513 1 3 7620 INVX1 $T=1595220 1410640 0 0 $X=1595218 $Y=1410238
X634 7519 1 3 7599 INVX1 $T=1603140 1158640 0 0 $X=1603138 $Y=1158238
X635 7558 1 3 7648 INVX1 $T=1605780 1360240 1 0 $X=1605778 $Y=1354800
X636 7553 1 3 7627 INVX1 $T=1605780 1390480 1 0 $X=1605778 $Y=1385040
X637 352 1 3 351 INVX1 $T=1609080 1219120 0 180 $X=1607760 $Y=1213680
X638 7329 1 3 7622 INVX1 $T=1608420 1319920 1 0 $X=1608418 $Y=1314480
X639 7544 1 3 7654 INVX1 $T=1611060 1340080 0 0 $X=1611058 $Y=1339678
X640 7708 1 3 7677 INVX1 $T=1625580 1269520 0 180 $X=1624260 $Y=1264080
X641 355 1 3 7396 INVX1 $T=1629540 1430800 1 0 $X=1629538 $Y=1425360
X642 7765 1 3 7800 INVX1 $T=1634820 1219120 1 0 $X=1634818 $Y=1213680
X643 7801 1 3 7839 INVX1 $T=1641420 1269520 0 180 $X=1640100 $Y=1264080
X644 7798 1 3 7786 INVX1 $T=1644720 1330000 0 180 $X=1643400 $Y=1324560
X645 7869 1 3 7876 INVX1 $T=1660560 1239280 1 0 $X=1660558 $Y=1233840
X646 7927 1 3 8015 INVX1 $T=1668480 1289680 0 0 $X=1668478 $Y=1289278
X647 7952 1 3 8035 INVX1 $T=1671120 1198960 1 0 $X=1671118 $Y=1193520
X648 8016 1 3 8041 INVX1 $T=1671120 1309840 0 0 $X=1671118 $Y=1309438
X649 7801 1 3 8166 INVX1 $T=1684320 1269520 1 0 $X=1684318 $Y=1264080
X650 8100 1 3 8147 INVX1 $T=1686960 1370320 1 0 $X=1686958 $Y=1364880
X651 363 1 3 370 INVX1 $T=1686960 1420720 1 0 $X=1686958 $Y=1415280
X652 7527 1 3 8247 INVX1 $T=1691580 1198960 0 0 $X=1691578 $Y=1198558
X653 7479 1 3 8188 INVX1 $T=1694880 1209040 0 0 $X=1694878 $Y=1208638
X654 8263 1 3 8240 INVX1 $T=1705440 1188880 1 0 $X=1705438 $Y=1183440
X655 8277 1 3 8244 INVX1 $T=1709400 1219120 0 180 $X=1708080 $Y=1213680
X656 8327 1 3 8251 INVX1 $T=1712040 1219120 1 180 $X=1710720 $Y=1218718
X657 8166 1 3 387 INVX1 $T=1715340 1239280 1 0 $X=1715338 $Y=1233840
X658 8335 1 3 8172 INVX1 $T=1717320 1198960 1 180 $X=1716000 $Y=1198558
X659 8477 1 3 8488 INVX1 $T=1741740 1289680 0 0 $X=1741738 $Y=1289278
X660 8633 1 3 8682 INVX1 $T=1765500 1209040 0 0 $X=1765498 $Y=1208638
X661 8658 1 3 8706 INVX1 $T=1770780 1198960 1 0 $X=1770778 $Y=1193520
X662 8729 1 3 8753 INVX1 $T=1782000 1239280 0 0 $X=1781998 $Y=1238878
X663 431 1 3 8750 INVX1 $T=1788600 1410640 1 0 $X=1788598 $Y=1405200
X664 8764 1 3 8883 INVX1 $T=1793880 1188880 0 0 $X=1793878 $Y=1188478
X665 8788 1 3 8704 INVX1 $T=1795200 1229200 0 180 $X=1793880 $Y=1223760
X666 8860 1 3 8807 INVX1 $T=1822920 1360240 0 0 $X=1822918 $Y=1359838
X667 410 1 3 9187 INVX1 $T=1844040 1430800 1 0 $X=1844038 $Y=1425360
X668 9235 1 3 9074 INVX1 $T=1851960 1168720 0 180 $X=1850640 $Y=1163280
X669 424 1 3 9188 INVX1 $T=1855260 1430800 1 0 $X=1855258 $Y=1425360
X670 9069 1 3 9323 INVX1 $T=1876380 1390480 0 0 $X=1876378 $Y=1390078
X671 9383 1 3 9353 INVX1 $T=1884300 1400560 1 180 $X=1882980 $Y=1400158
X672 9438 1 3 9359 INVX1 $T=1897500 1370320 1 180 $X=1896180 $Y=1369918
X673 9687 1 3 9756 INVX1 $T=1932480 1198960 0 0 $X=1932478 $Y=1198558
X674 9710 1 3 9780 INVX1 $T=1935120 1249360 1 0 $X=1935118 $Y=1243920
X675 9632 1 3 9766 INVX1 $T=1935120 1350160 1 0 $X=1935118 $Y=1344720
X676 435 1 3 9791 INVX1 $T=1937760 1219120 1 0 $X=1937758 $Y=1213680
X677 9386 1 3 9764 INVX1 $T=1937760 1249360 0 0 $X=1937758 $Y=1248958
X678 9736 1 3 9771 INVX1 $T=1943040 1209040 1 0 $X=1943038 $Y=1203600
X679 9735 1 3 9812 INVX1 $T=1948320 1229200 0 0 $X=1948318 $Y=1228798
X680 9508 1 3 9929 INVX1 $T=1969440 1239280 0 0 $X=1969438 $Y=1238878
X681 9792 1 3 9924 INVX1 $T=1976040 1340080 0 180 $X=1974720 $Y=1334640
X682 9684 1 3 9951 INVX1 $T=1978680 1319920 1 180 $X=1977360 $Y=1319518
X683 10148 1 3 10144 INVX1 $T=2013660 1420720 0 0 $X=2013658 $Y=1420318
X684 10318 1 3 10260 INVX1 $T=2025540 1219120 1 180 $X=2024220 $Y=1218718
X685 10264 1 3 10270 INVX1 $T=2028180 1299760 0 180 $X=2026860 $Y=1294320
X686 10325 1 3 10318 INVX1 $T=2033460 1229200 0 180 $X=2032140 $Y=1223760
X687 10396 1 3 10294 INVX1 $T=2046000 1148560 0 0 $X=2045998 $Y=1148158
X688 557 1 3 10316 INVX1 $T=2065140 1219120 1 180 $X=2063820 $Y=1218718
X689 560 1 3 10476 INVX1 $T=2067780 1269520 0 180 $X=2066460 $Y=1264080
X690 555 1 3 10497 INVX1 $T=2075040 1360240 1 180 $X=2073720 $Y=1359838
X691 549 1 3 10580 INVX1 $T=2090880 1340080 0 180 $X=2089560 $Y=1334640
X692 573 1 3 563 INVX1 $T=2104080 1178800 0 180 $X=2102760 $Y=1173360
X693 554 1 3 10701 INVX1 $T=2105400 1370320 1 0 $X=2105398 $Y=1364880
X694 579 1 3 584 INVX1 $T=2118600 1430800 1 0 $X=2118598 $Y=1425360
X695 558 1 3 10862 INVX1 $T=2126520 1330000 0 0 $X=2126518 $Y=1329598
X696 555 1 3 10941 INVX1 $T=2139060 1330000 1 180 $X=2137740 $Y=1329598
X697 549 1 3 10925 INVX1 $T=2140380 1309840 1 180 $X=2139060 $Y=1309438
X698 573 1 3 11091 INVX1 $T=2161500 1279600 0 180 $X=2160180 $Y=1274160
X699 11094 1 3 11180 INVX1 $T=2168100 1420720 1 0 $X=2168098 $Y=1415280
X700 553 1 3 568 INVX1 $T=2183940 1148560 1 0 $X=2183938 $Y=1143120
X701 560 1 3 11250 INVX1 $T=2188560 1350160 1 0 $X=2188558 $Y=1344720
X702 10172 1 3 11390 INVX1 $T=2211000 1219120 1 0 $X=2210998 $Y=1213680
X703 11449 1 3 11454 INVX1 $T=2217600 1360240 0 0 $X=2217598 $Y=1359838
X704 11445 1 3 11450 INVX1 $T=2220240 1370320 1 0 $X=2220238 $Y=1364880
X705 11254 1 3 610 INVX1 $T=2233440 1148560 1 0 $X=2233438 $Y=1143120
X706 551 1 3 11598 INVX1 $T=2238720 1158640 1 0 $X=2238718 $Y=1153200
X707 553 1 3 11538 INVX1 $T=2240040 1198960 1 180 $X=2238720 $Y=1198558
X708 559 1 3 11619 INVX1 $T=2250600 1178800 1 180 $X=2249280 $Y=1178398
X709 531 1 3 11814 INVX1 $T=2262480 1168720 0 0 $X=2262478 $Y=1168318
X710 615 1 3 11739 INVX1 $T=2267760 1410640 1 180 $X=2266440 $Y=1410238
X711 616 1 3 11738 INVX1 $T=2277000 1410640 0 180 $X=2275680 $Y=1405200
X712 609 1 3 11761 INVX1 $T=2277660 1138480 1 180 $X=2276340 $Y=1138078
X713 543 1 3 11736 INVX1 $T=2278320 1219120 0 0 $X=2278318 $Y=1218718
X714 11250 1 3 11883 INVX1 $T=2281620 1239280 0 0 $X=2281618 $Y=1238878
X715 573 1 3 11912 INVX1 $T=2288220 1239280 0 0 $X=2288218 $Y=1238878
X716 605 1 3 12042 INVX1 $T=2304060 1168720 0 0 $X=2304058 $Y=1168318
X717 11964 1 3 12070 INVX1 $T=2306700 1360240 0 0 $X=2306698 $Y=1359838
X718 12041 1 3 11937 INVX1 $T=2308020 1390480 0 180 $X=2306700 $Y=1385040
X719 12127 1 3 12292 INVX1 $T=2327160 1198960 1 0 $X=2327158 $Y=1193520
X720 12160 1 3 12271 INVX1 $T=2333100 1269520 0 0 $X=2333098 $Y=1269118
X721 12221 1 3 12275 INVX1 $T=2335080 1370320 1 0 $X=2335078 $Y=1364880
X722 12272 1 3 12437 INVX1 $T=2358840 1289680 0 0 $X=2358838 $Y=1289278
X723 12325 1 3 12462 INVX1 $T=2366760 1168720 1 0 $X=2366758 $Y=1163280
X724 12456 1 3 12465 INVX1 $T=2366760 1188880 0 0 $X=2366758 $Y=1188478
X725 12398 1 3 12463 INVX1 $T=2366760 1289680 1 0 $X=2366758 $Y=1284240
X726 12397 1 3 12402 INVX1 $T=2370720 1410640 1 180 $X=2369400 $Y=1410238
X727 12423 1 3 12496 INVX1 $T=2372040 1239280 1 0 $X=2372038 $Y=1233840
X728 12369 1 3 12495 INVX1 $T=2377320 1188880 0 0 $X=2377318 $Y=1188478
X729 12395 1 3 12527 INVX1 $T=2377320 1209040 0 0 $X=2377318 $Y=1208638
X730 12161 1 3 12622 INVX1 $T=2395800 1209040 0 0 $X=2395798 $Y=1208638
X731 12713 1 3 12427 INVX1 $T=2399100 1410640 0 180 $X=2397780 $Y=1405200
X732 12492 1 3 12714 INVX1 $T=2400420 1219120 0 0 $X=2400418 $Y=1218718
X733 12535 1 3 12715 INVX1 $T=2403720 1229200 1 0 $X=2403718 $Y=1223760
X734 12818 1 3 12868 INVX1 $T=2420880 1158640 0 0 $X=2420878 $Y=1158238
X735 637 1 3 12904 INVX1 $T=2426820 1148560 1 0 $X=2426818 $Y=1143120
X736 12874 1 3 12770 INVX1 $T=2428140 1410640 0 180 $X=2426820 $Y=1405200
X737 12906 1 3 12808 INVX1 $T=2433420 1390480 0 180 $X=2432100 $Y=1385040
X738 638 1 3 12909 INVX1 $T=2433420 1148560 1 0 $X=2433418 $Y=1143120
X739 12928 1 3 12929 INVX1 $T=2445300 1330000 1 0 $X=2445298 $Y=1324560
X740 643 1 3 13117 INVX1 $T=2447940 1410640 1 0 $X=2447938 $Y=1405200
X741 642 1 3 13088 INVX1 $T=2450580 1420720 0 0 $X=2450578 $Y=1420318
X742 13123 1 3 12888 INVX1 $T=2454540 1360240 0 180 $X=2453220 $Y=1354800
X743 13087 1 3 13089 INVX1 $T=2455860 1410640 0 0 $X=2455858 $Y=1410238
X744 13128 1 3 13278 INVX1 $T=2463780 1158640 0 0 $X=2463778 $Y=1158238
X745 13116 1 3 13001 INVX1 $T=2469060 1319920 1 0 $X=2469058 $Y=1314480
X746 13216 1 3 13239 INVX1 $T=2476980 1350160 1 0 $X=2476978 $Y=1344720
X747 647 1 3 13185 INVX1 $T=2483580 1400560 0 180 $X=2482260 $Y=1395120
X748 652 1 3 13282 INVX1 $T=2490180 1400560 0 180 $X=2488860 $Y=1395120
X749 13308 1 3 659 INVX1 $T=2494800 1410640 0 0 $X=2494798 $Y=1410238
X750 13335 1 3 13301 INVX1 $T=2497440 1269520 0 0 $X=2497438 $Y=1269118
X751 13424 1 3 13279 INVX1 $T=2501400 1188880 1 180 $X=2500080 $Y=1188478
X752 13420 1 3 13218 INVX1 $T=2502720 1370320 1 180 $X=2501400 $Y=1369918
X753 13287 1 3 13465 INVX1 $T=2514600 1188880 1 180 $X=2513280 $Y=1188478
X754 13500 1 3 13509 INVX1 $T=2513940 1340080 1 0 $X=2513938 $Y=1334640
X755 13519 1 3 13461 INVX1 $T=2515920 1370320 0 180 $X=2514600 $Y=1364880
X756 13680 1 3 13655 INVX1 $T=2533080 1340080 0 180 $X=2531760 $Y=1334640
X757 13679 1 3 13605 INVX1 $T=2533740 1309840 1 0 $X=2533738 $Y=1304400
X758 13610 1 3 13744 INVX1 $T=2539680 1309840 0 0 $X=2539678 $Y=1309438
X759 13743 1 3 13684 INVX1 $T=2541000 1410640 0 180 $X=2539680 $Y=1405200
X760 13787 1 3 13769 INVX1 $T=2546280 1340080 1 180 $X=2544960 $Y=1339678
X761 13874 1 3 13774 INVX1 $T=2551560 1178800 1 180 $X=2550240 $Y=1178398
X762 13875 1 3 13882 INVX1 $T=2553540 1340080 0 0 $X=2553538 $Y=1339678
X763 674 1 3 13938 INVX1 $T=2560140 1148560 0 0 $X=2560138 $Y=1148158
X764 676 1 3 679 INVX1 $T=2560800 1148560 1 0 $X=2560798 $Y=1143120
X765 13813 1 3 13833 INVX1 $T=2562120 1309840 1 180 $X=2560800 $Y=1309438
X766 13931 1 3 13912 INVX1 $T=2562120 1370320 1 180 $X=2560800 $Y=1369918
X767 13975 1 3 13899 INVX1 $T=2566740 1259440 1 180 $X=2565420 $Y=1259038
X768 13966 1 3 13834 INVX1 $T=2568060 1319920 1 180 $X=2566740 $Y=1319518
X769 13967 1 3 673 INVX1 $T=2570700 1309840 1 180 $X=2569380 $Y=1309438
X770 13808 1 3 13942 INVX1 $T=2570700 1269520 0 0 $X=2570698 $Y=1269118
X771 14011 1 3 13934 INVX1 $T=2572020 1239280 1 180 $X=2570700 $Y=1238878
X772 13876 1 3 13939 INVX1 $T=2574660 1259440 1 180 $X=2573340 $Y=1259038
X773 683 1 3 14009 INVX1 $T=2574000 1410640 0 0 $X=2573998 $Y=1410238
X774 13835 1 3 14035 INVX1 $T=2581260 1289680 1 0 $X=2581258 $Y=1284240
X775 14079 1 3 14020 INVX1 $T=2586540 1319920 0 0 $X=2586538 $Y=1319518
X776 14042 1 3 14111 INVX1 $T=2589180 1279600 0 0 $X=2589178 $Y=1279198
X777 14106 1 3 14227 INVX1 $T=2594460 1319920 1 0 $X=2594458 $Y=1314480
X778 14073 1 3 14232 INVX1 $T=2602380 1239280 0 0 $X=2602378 $Y=1238878
X779 14230 1 3 14115 INVX1 $T=2603700 1309840 0 180 $X=2602380 $Y=1304400
X780 14088 1 3 14310 INVX1 $T=2604360 1259440 0 0 $X=2604358 $Y=1259038
X781 14257 1 3 14311 INVX1 $T=2615580 1380400 1 0 $X=2615578 $Y=1374960
X782 14313 1 3 14279 INVX1 $T=2617560 1239280 1 180 $X=2616240 $Y=1238878
X783 14090 1 3 14338 INVX1 $T=2620860 1370320 0 0 $X=2620858 $Y=1369918
X784 14010 1 3 14277 INVX1 $T=2626140 1370320 0 0 $X=2626138 $Y=1369918
X785 1544 66 3 1543 1564 1 AOI21X2 $T=676500 1269520 0 180 $X=671880 $Y=1264080
X786 1600 66 3 1571 1596 1 AOI21X2 $T=681780 1239280 1 180 $X=677160 $Y=1238878
X787 1664 1870 3 1885 1886 1 AOI21X2 $T=721380 1259440 1 0 $X=721378 $Y=1254000
X788 1869 66 3 1889 1925 1 AOI21X2 $T=722700 1239280 1 0 $X=722698 $Y=1233840
X789 2767 2635 3 2761 2765 1 AOI21X2 $T=853380 1178800 1 180 $X=848760 $Y=1178398
X790 2868 2843 3 2767 2872 1 AOI21X2 $T=873840 1178800 1 0 $X=873838 $Y=1173360
X791 117 3020 3 3059 3067 1 AOI21X2 $T=898920 1148560 1 0 $X=898918 $Y=1143120
X792 3137 3142 3 3160 120 1 AOI21X2 $T=920700 1158640 1 0 $X=920698 $Y=1153200
X793 3403 3378 3 3412 3374 1 AOI21X2 $T=959640 1299760 1 0 $X=959638 $Y=1294320
X794 3732 3738 3 3749 3695 1 AOI21X2 $T=1011780 1259440 1 0 $X=1011778 $Y=1254000
X795 3745 3749 3 3744 3771 1 AOI21X2 $T=1016400 1229200 0 180 $X=1011780 $Y=1223760
X796 3861 3856 3 3900 3778 1 AOI21X2 $T=1035540 1360240 0 0 $X=1035538 $Y=1359838
X797 6405 6402 3 6428 6437 1 AOI21X2 $T=1430220 1188880 1 0 $X=1430218 $Y=1183440
X798 6458 6457 3 6566 6658 1 AOI21X2 $T=1447380 1279600 0 0 $X=1447378 $Y=1279198
X799 6759 6841 3 6847 6827 1 AOI21X2 $T=1492920 1330000 0 0 $X=1492918 $Y=1329598
X800 6737 6790 3 6836 6921 1 AOI21X2 $T=1494240 1158640 1 0 $X=1494238 $Y=1153200
X801 6947 6702 3 6790 6879 1 AOI21X2 $T=1505460 1168720 1 180 $X=1500840 $Y=1168318
X802 6978 7031 3 7088 7072 1 AOI21X2 $T=1529880 1219120 0 0 $X=1529878 $Y=1218718
X803 7179 7127 3 7031 7166 1 AOI21X2 $T=1544400 1239280 1 180 $X=1539780 $Y=1238878
X804 7260 7103 3 7257 7278 1 AOI21X2 $T=1557600 1350160 1 180 $X=1552980 $Y=1349758
X805 7837 7875 3 7800 7917 1 AOI21X2 $T=1651980 1219120 0 180 $X=1647360 $Y=1213680
X806 8731 8682 3 8706 8728 1 AOI21X2 $T=1782660 1198960 1 180 $X=1778040 $Y=1198558
X807 8749 8755 3 8753 8788 1 AOI21X2 $T=1789260 1239280 0 0 $X=1789258 $Y=1238878
X808 10319 10260 3 10377 545 1 AOI21X2 $T=2045340 1178800 0 180 $X=2040720 $Y=1173360
X809 547 10294 3 10384 546 1 AOI21X2 $T=2046660 1148560 0 180 $X=2042040 $Y=1143120
X810 11451 11454 3 11450 11303 1 AOI21X2 $T=2219580 1370320 1 180 $X=2214960 $Y=1369918
X811 11451 11581 3 11444 11578 1 AOI21X2 $T=2240700 1350160 1 180 $X=2236080 $Y=1349758
X812 11586 11444 3 11599 11620 1 AOI21X2 $T=2244660 1330000 0 180 $X=2240040 $Y=1324560
X813 11734 11738 3 11739 11703 1 AOI21X2 $T=2256540 1410640 1 0 $X=2256538 $Y=1405200
X814 11734 11847 3 11849 11844 1 AOI21X2 $T=2275020 1390480 0 0 $X=2275018 $Y=1390078
X815 618 12328 3 626 12244 1 AOI21X2 $T=2350920 1420720 0 180 $X=2346300 $Y=1415280
X816 618 12323 3 12327 12320 1 AOI21X2 $T=2346960 1410640 0 0 $X=2346958 $Y=1410238
X817 626 12503 3 12536 12537 1 AOI21X2 $T=2377320 1410640 1 0 $X=2377318 $Y=1405200
X818 12999 12929 3 13001 13039 1 AOI21X2 $T=2445960 1319920 1 0 $X=2445958 $Y=1314480
X819 13099 13117 3 13179 13219 1 AOI21X2 $T=2469060 1410640 1 0 $X=2469058 $Y=1405200
X820 13222 13317 3 13339 13269 1 AOI21X2 $T=2494800 1198960 0 0 $X=2494798 $Y=1198558
X821 13589 13339 3 13691 13597 1 AOI21X2 $T=2531100 1188880 0 0 $X=2531098 $Y=1188478
X822 13744 13814 3 13833 13808 1 AOI21X2 $T=2546940 1309840 0 0 $X=2546938 $Y=1309438
X823 3 1545 58 1567 1 NOR2X1 $T=670560 1289680 0 180 $X=668580 $Y=1284240
X824 3 58 62 1544 1 NOR2X1 $T=669240 1259440 0 0 $X=669238 $Y=1259038
X825 3 64 1541 1574 1 NOR2X1 $T=671220 1209040 1 0 $X=671218 $Y=1203600
X826 3 1574 1605 1597 1 NOR2X1 $T=682440 1219120 0 0 $X=682438 $Y=1218718
X827 3 1752 1672 1636 1 NOR2X1 $T=696960 1350160 1 180 $X=694980 $Y=1349758
X828 3 1840 62 1869 1 NOR2X1 $T=718740 1239280 0 0 $X=718738 $Y=1238878
X829 3 79 1865 1839 1 NOR2X1 $T=720720 1289680 0 0 $X=720718 $Y=1289278
X830 3 1996 1918 2012 1 NOR2X1 $T=742500 1420720 0 0 $X=742498 $Y=1420318
X831 3 2113 2047 1782 1 NOR2X1 $T=749760 1370320 1 180 $X=747780 $Y=1369918
X832 3 88 86 1918 1 NOR2X1 $T=752400 1430800 0 180 $X=750420 $Y=1425360
X833 3 2142 2166 2108 1 NOR2X1 $T=761640 1350160 1 180 $X=759660 $Y=1349758
X834 3 89 2182 1996 1 NOR2X1 $T=766260 1420720 0 180 $X=764280 $Y=1415280
X835 3 2236 2232 2142 1 NOR2X1 $T=771540 1340080 1 180 $X=769560 $Y=1339678
X836 3 2215 2237 2212 1 NOR2X1 $T=770880 1269520 0 0 $X=770878 $Y=1269118
X837 3 2309 2242 2215 1 NOR2X1 $T=774180 1299760 1 180 $X=772200 $Y=1299358
X838 3 2208 2245 2047 1 NOR2X1 $T=774840 1390480 0 180 $X=772860 $Y=1385040
X839 3 2307 2282 2113 1 NOR2X1 $T=780780 1370320 1 180 $X=778800 $Y=1369918
X840 3 2313 2302 2271 1 NOR2X1 $T=783420 1188880 1 180 $X=781440 $Y=1188478
X841 3 91 2269 2214 1 NOR2X1 $T=786060 1168720 0 180 $X=784080 $Y=1163280
X842 3 2342 2336 2166 1 NOR2X1 $T=787380 1350160 1 180 $X=785400 $Y=1349758
X843 3 2404 2371 2281 1 NOR2X1 $T=792660 1279600 1 180 $X=790680 $Y=1279198
X844 3 2403 2380 2313 1 NOR2X1 $T=799260 1188880 1 180 $X=797280 $Y=1188478
X845 3 2543 2518 2321 1 NOR2X1 $T=817740 1279600 0 180 $X=815760 $Y=1274160
X846 3 115 2869 2844 1 NOR2X1 $T=871200 1219120 0 180 $X=869220 $Y=1213680
X847 3 3119 3184 3192 1 NOR2X1 $T=927960 1400560 0 0 $X=927958 $Y=1400158
X848 3 3404 3357 3373 1 NOR2X1 $T=958980 1239280 1 180 $X=957000 $Y=1238878
X849 3 3434 3416 3248 1 NOR2X1 $T=964260 1309840 0 180 $X=962280 $Y=1304400
X850 3 141 140 3404 1 NOR2X1 $T=976140 1239280 1 180 $X=974160 $Y=1238878
X851 3 3694 3671 143 1 NOR2X1 $T=1004520 1168720 0 180 $X=1002540 $Y=1163280
X852 3 3812 3704 3736 1 NOR2X1 $T=1013100 1330000 0 180 $X=1011120 $Y=1324560
X853 3 3707 3793 3745 1 NOR2X1 $T=1019040 1239280 1 0 $X=1019038 $Y=1233840
X854 3 3841 3796 3671 1 NOR2X1 $T=1030920 1188880 0 180 $X=1028940 $Y=1183440
X855 3 4031 3903 3803 1 NOR2X1 $T=1040820 1259440 1 180 $X=1038840 $Y=1259038
X856 3 3924 3803 3738 1 NOR2X1 $T=1040820 1269520 0 180 $X=1038840 $Y=1264080
X857 3 3906 3877 3704 1 NOR2X1 $T=1040160 1330000 0 0 $X=1040158 $Y=1329598
X858 3 4266 4146 4120 1 NOR2X1 $T=1080420 1390480 1 180 $X=1078440 $Y=1390078
X859 3 191 4459 4666 1 NOR2X1 $T=1162920 1209040 1 180 $X=1160940 $Y=1208638
X860 3 232 191 4990 1 NOR2X1 $T=1209780 1279600 0 180 $X=1207800 $Y=1274160
X861 3 230 199 5022 1 NOR2X1 $T=1222320 1229200 0 0 $X=1222318 $Y=1228798
X862 3 5463 5191 5542 1 NOR2X1 $T=1286340 1209040 1 0 $X=1286338 $Y=1203600
X863 3 186 6105 6099 1 NOR2X1 $T=1386000 1340080 0 0 $X=1385998 $Y=1339678
X864 3 5614 6087 6280 1 NOR2X1 $T=1396560 1289680 1 0 $X=1396558 $Y=1284240
X865 3 6044 6253 6282 1 NOR2X1 $T=1401180 1249360 1 0 $X=1401178 $Y=1243920
X866 3 6282 6307 6341 1 NOR2X1 $T=1409100 1239280 0 0 $X=1409098 $Y=1238878
X867 3 5649 6595 6598 1 NOR2X1 $T=1455300 1249360 0 0 $X=1455298 $Y=1248958
X868 3 320 3093 6694 1 NOR2X1 $T=1469160 1299760 0 180 $X=1467180 $Y=1294320
X869 3 6806 6821 323 1 NOR2X1 $T=1490280 1420720 0 0 $X=1490278 $Y=1420318
X870 3 331 6998 7032 1 NOR2X1 $T=1525260 1279600 1 0 $X=1525258 $Y=1274160
X871 3 331 334 7129 1 NOR2X1 $T=1537800 1299760 1 0 $X=1537798 $Y=1294320
X872 3 7138 6998 7161 1 NOR2X1 $T=1542420 1279600 1 0 $X=1542418 $Y=1274160
X873 3 3246 7284 7287 1 NOR2X1 $T=1557600 1209040 1 0 $X=1557598 $Y=1203600
X874 3 340 7376 339 1 NOR2X1 $T=1571460 1138480 0 0 $X=1571458 $Y=1138078
X875 3 342 338 7406 1 NOR2X1 $T=1581360 1259440 1 180 $X=1579380 $Y=1259038
X876 3 7283 7384 7383 1 NOR2X1 $T=1582020 1239280 1 0 $X=1582018 $Y=1233840
X877 3 363 362 360 1 NOR2X1 $T=1654620 1410640 1 180 $X=1652640 $Y=1410238
X878 3 370 367 365 1 NOR2X1 $T=1667820 1420720 0 180 $X=1665840 $Y=1415280
X879 3 8173 6666 8270 1 NOR2X1 $T=1704780 1350160 1 0 $X=1704778 $Y=1344720
X880 3 8628 6852 8590 1 NOR2X1 $T=1760880 1269520 0 180 $X=1758900 $Y=1264080
X881 3 356 440 8884 1 NOR2X1 $T=1795860 1410640 1 0 $X=1795858 $Y=1405200
X882 3 8887 8882 8784 1 NOR2X1 $T=1807080 1158640 0 180 $X=1805100 $Y=1153200
X883 3 10268 535 10148 1 NOR2X1 $T=2016960 1420720 1 180 $X=2014980 $Y=1420318
X884 3 10302 10299 10298 1 NOR2X1 $T=2030160 1239280 0 180 $X=2028180 $Y=1233840
X885 3 10316 10297 10323 1 NOR2X1 $T=2032140 1209040 1 0 $X=2032138 $Y=1203600
X886 3 10356 10323 10319 1 NOR2X1 $T=2034120 1178800 0 180 $X=2032140 $Y=1173360
X887 3 10238 10266 10356 1 NOR2X1 $T=2046660 1188880 1 0 $X=2046658 $Y=1183440
X888 3 10520 10531 10530 1 NOR2X1 $T=2074380 1279600 0 180 $X=2072400 $Y=1274160
X889 3 10623 10633 569 1 NOR2X1 $T=2086260 1410640 1 0 $X=2086258 $Y=1405200
X890 3 10648 10621 10629 1 NOR2X1 $T=2094180 1319920 1 180 $X=2092200 $Y=1319518
X891 3 10572 10580 10621 1 NOR2X1 $T=2094180 1330000 1 180 $X=2092200 $Y=1329598
X892 3 10558 562 10648 1 NOR2X1 $T=2096160 1319920 1 0 $X=2096158 $Y=1314480
X893 3 10702 10823 10784 1 NOR2X1 $T=2115300 1370320 1 0 $X=2115298 $Y=1364880
X894 3 10860 10784 10863 1 NOR2X1 $T=2120580 1400560 0 0 $X=2120578 $Y=1400158
X895 3 10866 10865 10860 1 NOR2X1 $T=2122560 1360240 0 180 $X=2120580 $Y=1354800
X896 3 587 593 598 1 NOR2X1 $T=2154900 1430800 1 0 $X=2154898 $Y=1425360
X897 3 11251 11232 11276 1 NOR2X1 $T=2197140 1410640 1 180 $X=2195160 $Y=1410238
X898 3 11125 11259 11251 1 NOR2X1 $T=2195820 1400560 1 0 $X=2195818 $Y=1395120
X899 3 11182 11357 11417 1 NOR2X1 $T=2209020 1340080 1 0 $X=2209018 $Y=1334640
X900 3 11285 11412 11449 1 NOR2X1 $T=2211000 1350160 0 0 $X=2210998 $Y=1349758
X901 3 11356 11512 11546 1 NOR2X1 $T=2229480 1319920 1 0 $X=2229478 $Y=1314480
X902 3 11449 11417 11581 1 NOR2X1 $T=2230140 1350160 1 0 $X=2230138 $Y=1344720
X903 3 11905 12072 12130 1 NOR2X1 $T=2308020 1148560 1 0 $X=2308018 $Y=1143120
X904 3 12102 11821 12161 1 NOR2X1 $T=2315940 1209040 0 180 $X=2313960 $Y=1203600
X905 3 621 11965 12270 1 NOR2X1 $T=2331120 1138480 0 0 $X=2331118 $Y=1138078
X906 3 11963 11962 12423 1 NOR2X1 $T=2344980 1229200 1 0 $X=2344978 $Y=1223760
X907 3 12220 12131 12369 1 NOR2X1 $T=2348940 1198960 1 0 $X=2348938 $Y=1193520
X908 3 12270 12130 629 1 NOR2X1 $T=2358840 1148560 1 0 $X=2358838 $Y=1143120
X909 3 12399 12221 12373 1 NOR2X1 $T=2361480 1360240 0 0 $X=2361478 $Y=1359838
X910 3 12435 12427 12397 1 NOR2X1 $T=2365440 1410640 0 180 $X=2363460 $Y=1405200
X911 3 12161 12466 12467 1 NOR2X1 $T=2368080 1209040 1 0 $X=2368078 $Y=1203600
X912 3 12522 12535 12565 1 NOR2X1 $T=2384580 1229200 1 0 $X=2384578 $Y=1223760
X913 3 12161 12714 12807 1 NOR2X1 $T=2400420 1219120 1 0 $X=2400418 $Y=1213680
X914 3 12534 12714 12746 1 NOR2X1 $T=2403720 1209040 0 0 $X=2403718 $Y=1208638
X915 3 12628 12808 12717 1 NOR2X1 $T=2418240 1370320 1 180 $X=2416260 $Y=1369918
X916 3 648 642 13099 1 NOR2X1 $T=2457840 1430800 1 0 $X=2457838 $Y=1425360
X917 3 653 645 654 1 NOR2X1 $T=2488200 1420720 0 0 $X=2488198 $Y=1420318
X918 3 13093 13655 13679 1 NOR2X1 $T=2529780 1319920 1 0 $X=2529778 $Y=1314480
X919 3 669 667 13743 1 NOR2X1 $T=2538360 1420720 0 0 $X=2538358 $Y=1420318
X920 3 13122 13769 13812 1 NOR2X1 $T=2545620 1158640 1 0 $X=2545618 $Y=1153200
X921 3 676 13812 13902 1 NOR2X1 $T=2552220 1158640 0 0 $X=2552218 $Y=1158238
X922 3 680 13900 13971 1 NOR2X1 $T=2568060 1380400 0 0 $X=2568058 $Y=1379998
X923 3 13835 14060 14089 1 NOR2X1 $T=2581260 1279600 1 0 $X=2581258 $Y=1274160
X924 3 14011 13975 14012 1 NOR2X1 $T=2583240 1259440 1 180 $X=2581260 $Y=1259038
X925 3 14071 14064 13985 1 NOR2X1 $T=2584560 1168720 0 180 $X=2582580 $Y=1163280
X926 3 14018 13898 14090 1 NOR2X1 $T=2586540 1410640 1 0 $X=2586538 $Y=1405200
X927 3 690 14115 14071 1 NOR2X1 $T=2592480 1178800 0 180 $X=2590500 $Y=1173360
X928 3 14110 691 14228 1 NOR2X1 $T=2593140 1350160 0 0 $X=2593138 $Y=1349758
X929 3 694 14227 14064 1 NOR2X1 $T=2608980 1158640 0 0 $X=2608978 $Y=1158238
X930 3 13876 14310 14309 1 NOR2X1 $T=2616900 1259440 0 0 $X=2616898 $Y=1259038
X931 61 45 1 3 1508 NOR2X2 $T=663960 1380400 0 0 $X=663958 $Y=1379998
X932 1601 68 1 3 1605 NOR2X2 $T=680460 1229200 0 0 $X=680458 $Y=1228798
X933 1839 1806 1 3 1549 NOR2X2 $T=712140 1279600 0 180 $X=708840 $Y=1274160
X934 1897 81 1 3 1806 NOR2X2 $T=735900 1279600 1 0 $X=735898 $Y=1274160
X935 2870 2841 1 3 2819 NOR2X2 $T=865260 1269520 0 180 $X=861960 $Y=1264080
X936 2689 2844 1 3 2843 NOR2X2 $T=871860 1198960 1 180 $X=868560 $Y=1198558
X937 2917 1812 1 3 2898 NOR2X2 $T=881760 1309840 1 180 $X=878460 $Y=1309438
X938 2942 3087 1 3 3060 NOR2X2 $T=910800 1340080 1 180 $X=907500 $Y=1339678
X939 2956 3119 1 3 3070 NOR2X2 $T=916080 1400560 1 180 $X=912780 $Y=1400158
X940 3114 122 1 3 3119 NOR2X2 $T=914100 1410640 0 0 $X=914098 $Y=1410238
X941 135 133 1 3 3357 NOR2X2 $T=960300 1249360 1 0 $X=960298 $Y=1243920
X942 3434 3475 1 3 3403 NOR2X2 $T=976800 1299760 1 0 $X=976798 $Y=1294320
X943 3557 146 1 3 3416 NOR2X2 $T=990000 1299760 1 0 $X=989998 $Y=1294320
X944 148 149 1 3 3434 NOR2X2 $T=995940 1309840 0 180 $X=992640 $Y=1304400
X945 151 154 1 3 3495 NOR2X2 $T=997260 1380400 0 180 $X=993960 $Y=1374960
X946 144 145 1 3 3475 NOR2X2 $T=995280 1299760 1 0 $X=995278 $Y=1294320
X947 3875 3902 1 3 3707 NOR2X2 $T=1027620 1249360 0 180 $X=1024320 $Y=1243920
X948 3904 3921 1 3 3694 NOR2X2 $T=1040160 1168720 0 180 $X=1036860 $Y=1163280
X949 3957 4022 1 3 3812 NOR2X2 $T=1043460 1319920 1 180 $X=1040160 $Y=1319518
X950 3905 3922 1 3 3793 NOR2X2 $T=1046100 1229200 0 0 $X=1046098 $Y=1228798
X951 4032 4027 1 3 3924 NOR2X2 $T=1052040 1279600 1 180 $X=1048740 $Y=1279198
X952 247 198 1 3 4778 NOR2X2 $T=1234860 1148560 0 0 $X=1234858 $Y=1148158
X953 6251 6149 1 3 6307 NOR2X2 $T=1401840 1229200 0 0 $X=1401838 $Y=1228798
X954 3224 310 1 3 6459 NOR2X2 $T=1439460 1420720 1 180 $X=1436160 $Y=1420318
X955 6339 6459 1 3 6481 NOR2X2 $T=1441440 1410640 1 0 $X=1441438 $Y=1405200
X956 3350 317 1 3 6485 NOR2X2 $T=1446720 1380400 0 180 $X=1443420 $Y=1374960
X957 6570 6006 1 3 6635 NOR2X2 $T=1450680 1219120 0 0 $X=1450678 $Y=1218718
X958 6627 6005 1 3 6664 NOR2X2 $T=1461240 1209040 0 0 $X=1461238 $Y=1208638
X959 3274 6696 1 3 6699 NOR2X2 $T=1467180 1269520 1 180 $X=1463880 $Y=1269118
X960 6699 6694 1 3 6727 NOR2X2 $T=1471140 1289680 1 0 $X=1471138 $Y=1284240
X961 6664 6635 1 3 6773 NOR2X2 $T=1487640 1219120 0 180 $X=1484340 $Y=1213680
X962 6977 6841 1 3 7001 NOR2X2 $T=1512060 1340080 1 0 $X=1512058 $Y=1334640
X963 7256 7011 1 3 7261 NOR2X2 $T=1552980 1370320 0 0 $X=1552978 $Y=1369918
X964 7321 7324 1 3 7320 NOR2X2 $T=1560900 1340080 0 0 $X=1560898 $Y=1339678
X965 7393 7180 1 3 7324 NOR2X2 $T=1572120 1330000 1 180 $X=1568820 $Y=1329598
X966 7519 7542 1 3 7547 NOR2X2 $T=1601160 1148560 1 180 $X=1597860 $Y=1148158
X967 7598 7626 1 3 7658 NOR2X2 $T=1618980 1239280 0 180 $X=1615680 $Y=1233840
X968 7932 7952 1 3 7986 NOR2X2 $T=1669140 1168720 0 0 $X=1669138 $Y=1168318
X969 8271 8246 1 3 8375 NOR2X2 $T=1733160 1390480 0 0 $X=1733158 $Y=1390078
X970 443 445 1 3 8860 NOR2X2 $T=1803120 1360240 0 180 $X=1799820 $Y=1354800
X971 7264 8919 1 3 8882 NOR2X2 $T=1809720 1138480 1 180 $X=1806420 $Y=1138078
X972 7009 8941 1 3 8887 NOR2X2 $T=1816320 1158640 0 180 $X=1813020 $Y=1153200
X973 473 474 1 3 9208 NOR2X2 $T=1861860 1148560 0 0 $X=1861858 $Y=1148158
X974 475 476 1 3 9121 NOR2X2 $T=1865160 1158640 1 180 $X=1861860 $Y=1158238
X975 9208 9121 1 3 9314 NOR2X2 $T=1865160 1158640 1 0 $X=1865158 $Y=1153200
X976 515 513 1 3 9732 NOR2X2 $T=1956240 1330000 1 180 $X=1952940 $Y=1329598
X977 544 542 1 3 10349 NOR2X2 $T=2035440 1330000 0 0 $X=2035438 $Y=1329598
X978 11553 11387 1 3 11585 NOR2X2 $T=2238060 1289680 0 0 $X=2238058 $Y=1289278
X979 11546 11585 1 3 11586 NOR2X2 $T=2242680 1319920 0 180 $X=2239380 $Y=1314480
X980 11927 11615 1 3 11960 NOR2X2 $T=2292840 1299760 0 0 $X=2292838 $Y=1299358
X981 12159 11805 1 3 12160 NOR2X2 $T=2321220 1269520 1 0 $X=2321218 $Y=1264080
X982 11811 11791 1 3 12274 NOR2X2 $T=2329140 1299760 1 0 $X=2329138 $Y=1294320
X983 12165 11827 1 3 12246 NOR2X2 $T=2337060 1249360 0 0 $X=2337058 $Y=1248958
X984 11926 11826 1 3 12396 NOR2X2 $T=2338380 1209040 0 0 $X=2338378 $Y=1208638
X985 12160 12246 1 3 12247 NOR2X2 $T=2341680 1269520 0 180 $X=2338380 $Y=1264080
X986 624 625 1 3 12328 NOR2X2 $T=2347620 1430800 1 0 $X=2347618 $Y=1425360
X987 11960 12274 1 3 12398 NOR2X2 $T=2355540 1299760 1 0 $X=2355538 $Y=1294320
X988 630 12434 1 3 12221 NOR2X2 $T=2362800 1370320 0 180 $X=2359500 $Y=1364880
X989 12423 12396 1 3 12492 NOR2X2 $T=2360820 1229200 1 0 $X=2360818 $Y=1223760
X990 12477 12397 1 3 12503 NOR2X2 $T=2370060 1410640 1 0 $X=2370058 $Y=1405200
X991 12770 12569 1 3 12477 NOR2X2 $T=2408340 1390480 0 0 $X=2408338 $Y=1390078
X992 12777 12717 1 3 12811 NOR2X2 $T=2410320 1370320 1 0 $X=2410318 $Y=1364880
X993 12888 12650 1 3 12777 NOR2X2 $T=2428800 1360240 1 0 $X=2428798 $Y=1354800
X994 656 13319 1 3 13306 NOR2X2 $T=2495460 1299760 1 180 $X=2492160 $Y=1299358
X995 13224 13318 1 3 13334 NOR2X2 $T=2497440 1249360 0 0 $X=2497438 $Y=1248958
X996 13427 13432 1 3 13430 NOR2X2 $T=2506020 1178800 0 0 $X=2506018 $Y=1178398
X997 13645 13609 1 3 13317 NOR2X2 $T=2529120 1219120 1 0 $X=2529118 $Y=1213680
X998 13287 13785 1 3 13589 NOR2X2 $T=2543640 1198960 0 180 $X=2540340 $Y=1193520
X999 13834 12722 1 3 13975 NOR2X2 $T=2567400 1259440 1 0 $X=2567398 $Y=1254000
X1000 14020 684 1 3 14011 NOR2X2 $T=2580600 1239280 0 0 $X=2580598 $Y=1238878
X1001 14073 14011 1 3 14088 NOR2X2 $T=2583240 1249360 0 0 $X=2583238 $Y=1248958
X1002 14309 14283 1 3 14224 NOR2X2 $T=2614260 1269520 1 0 $X=2614258 $Y=1264080
X1003 108 99 1 3 2399 OR2XL $T=825660 1209040 1 180 $X=823020 $Y=1208638
X1004 87 97 1 3 2567 OR2XL $T=826980 1380400 0 180 $X=824340 $Y=1374960
X1005 108 110 1 3 2521 OR2XL $T=829620 1299760 1 180 $X=826980 $Y=1299358
X1006 99 106 1 3 2517 OR2XL $T=829620 1390480 1 180 $X=826980 $Y=1390078
X1007 2875 56 1 3 2922 OR2XL $T=879120 1259440 0 0 $X=879118 $Y=1259038
X1008 184 185 1 3 4360 OR2XL $T=1098900 1309840 1 0 $X=1098898 $Y=1304400
X1009 184 4615 1 3 4617 OR2XL $T=1152360 1360240 0 0 $X=1152358 $Y=1359838
X1010 187 242 1 3 5103 OR2XL $T=1213080 1410640 0 0 $X=1213078 $Y=1410238
X1011 5489 5433 1 3 5652 OR2XL $T=1288980 1158640 1 0 $X=1288978 $Y=1153200
X1012 138 5849 1 3 5944 OR2XL $T=1346400 1410640 1 0 $X=1346398 $Y=1405200
X1013 136 6028 1 3 5998 OR2XL $T=1372140 1390480 0 180 $X=1369500 $Y=1385040
X1014 298 6028 1 3 6001 OR2XL $T=1370820 1380400 1 0 $X=1370818 $Y=1374960
X1015 179 6123 1 3 6190 OR2XL $T=1386660 1390480 1 0 $X=1386658 $Y=1385040
X1016 6342 8152 1 3 8154 OR2XL $T=1692900 1360240 1 0 $X=1692898 $Y=1354800
X1017 470 9188 1 3 9204 OR2XL $T=1851300 1430800 1 0 $X=1851298 $Y=1425360
X1018 633 12502 1 3 12457 OR2XL $T=2377980 1350160 0 180 $X=2375340 $Y=1344720
X1019 12042 609 1 3 12835 OR2XL $T=2409660 1158640 0 0 $X=2409658 $Y=1158238
X1020 2875 56 2937 1 3 NAND2X2 $T=879780 1249360 1 180 $X=876480 $Y=1248958
X1021 2917 1812 2948 1 3 NAND2X2 $T=882420 1319920 0 180 $X=879120 $Y=1314480
X1022 2939 60 2984 1 3 NAND2X2 $T=887040 1350160 1 0 $X=887038 $Y=1344720
X1023 2941 2842 2953 1 3 NAND2X2 $T=892320 1209040 0 0 $X=892318 $Y=1208638
X1024 2951 116 3015 1 3 NAND2X2 $T=894960 1370320 0 0 $X=894958 $Y=1369918
X1025 3064 59 3022 1 3 NAND2X2 $T=899580 1330000 1 180 $X=896280 $Y=1329598
X1026 3114 122 3134 1 3 NAND2X2 $T=914760 1420720 0 180 $X=911460 $Y=1415280
X1027 3408 127 3436 1 3 NAND2X2 $T=961620 1410640 1 0 $X=961618 $Y=1405200
X1028 135 133 3273 1 3 NAND2X2 $T=972180 1249360 1 0 $X=972178 $Y=1243920
X1029 151 154 3481 1 3 NAND2X2 $T=1001880 1380400 1 0 $X=1001878 $Y=1374960
X1030 3745 3738 3735 1 3 NAND2X2 $T=1012440 1239280 1 0 $X=1012438 $Y=1233840
X1031 4032 4027 3801 1 3 NAND2X2 $T=1054680 1289680 1 0 $X=1054678 $Y=1284240
X1032 201 4438 4435 1 3 NAND2X2 $T=1122000 1420720 1 180 $X=1118700 $Y=1420318
X1033 226 4726 4753 1 3 NAND2X2 $T=1179420 1420720 0 180 $X=1176120 $Y=1415280
X1034 251 5110 5188 1 3 NAND2X2 $T=1232220 1420720 0 0 $X=1232218 $Y=1420318
X1035 3224 310 6434 1 3 NAND2X2 $T=1439460 1410640 1 180 $X=1436160 $Y=1410238
X1036 315 3423 6593 1 3 NAND2X2 $T=1452000 1360240 0 0 $X=1451998 $Y=1359838
X1037 317 3350 6630 1 3 NAND2X2 $T=1454640 1380400 1 0 $X=1454638 $Y=1374960
X1038 6570 6006 6575 1 3 NAND2X2 $T=1457940 1229200 0 180 $X=1454640 $Y=1223760
X1039 6629 5994 6792 1 3 NAND2X2 $T=1474440 1178800 1 180 $X=1471140 $Y=1178398
X1040 320 3093 6753 1 3 NAND2X2 $T=1477080 1309840 1 0 $X=1477078 $Y=1304400
X1041 3355 7005 7027 1 3 NAND2X2 $T=1524600 1249360 0 180 $X=1521300 $Y=1243920
X1042 7055 6920 7092 1 3 NAND2X2 $T=1527240 1390480 1 0 $X=1527238 $Y=1385040
X1043 7256 7011 7214 1 3 NAND2X2 $T=1552980 1370320 1 180 $X=1549680 $Y=1369918
X1044 2944 7176 7255 1 3 NAND2X2 $T=1554300 1178800 0 180 $X=1551000 $Y=1173360
X1045 3246 7284 7378 1 3 NAND2X2 $T=1567500 1209040 0 180 $X=1564200 $Y=1203600
X1046 2820 7391 7377 1 3 NAND2X2 $T=1574100 1158640 0 180 $X=1570800 $Y=1153200
X1047 7418 7378 7443 1 3 NAND2X2 $T=1578720 1198960 0 0 $X=1578718 $Y=1198558
X1048 7478 7285 7542 1 3 NAND2X2 $T=1591920 1178800 0 0 $X=1591918 $Y=1178398
X1049 7392 7604 7602 1 3 NAND2X2 $T=1608420 1299760 1 180 $X=1605120 $Y=1299358
X1050 7258 7597 7625 1 3 NAND2X2 $T=1611060 1249360 0 180 $X=1607760 $Y=1243920
X1051 7764 7837 7960 1 3 NAND2X2 $T=1651980 1219120 0 0 $X=1651978 $Y=1218718
X1052 7836 7982 7981 1 3 NAND2X2 $T=1664520 1168720 1 180 $X=1661220 $Y=1168318
X1053 8151 379 8144 1 3 NAND2X2 $T=1694220 1158640 1 180 $X=1690920 $Y=1158238
X1054 378 8295 8148 1 3 NAND2X2 $T=1694880 1148560 1 180 $X=1691580 $Y=1148158
X1055 8731 8653 8785 1 3 NAND2X2 $T=1781340 1209040 1 0 $X=1781338 $Y=1203600
X1056 443 445 8861 1 3 NAND2X2 $T=1803120 1350160 1 180 $X=1799820 $Y=1349758
X1057 7009 8941 8892 1 3 NAND2X2 $T=1815660 1168720 0 180 $X=1812360 $Y=1163280
X1058 9537 9536 9399 1 3 NAND2X2 $T=1906740 1309840 1 0 $X=1906738 $Y=1304400
X1059 9689 9665 9684 1 3 NAND2X2 $T=1932480 1340080 1 180 $X=1929180 $Y=1339678
X1060 9883 9868 9708 1 3 NAND2X2 $T=1959540 1299760 1 0 $X=1959538 $Y=1294320
X1061 530 529 10051 1 3 NAND2X2 $T=1997820 1249360 0 0 $X=1997818 $Y=1248958
X1062 536 537 10170 1 3 NAND2X2 $T=2018280 1269520 0 0 $X=2018278 $Y=1269118
X1063 539 540 10272 1 3 NAND2X2 $T=2030160 1309840 1 0 $X=2030158 $Y=1304400
X1064 542 544 10295 1 3 NAND2X2 $T=2034780 1340080 1 0 $X=2034778 $Y=1334640
X1065 11586 11581 11596 1 3 NAND2X2 $T=2242680 1340080 0 180 $X=2239380 $Y=1334640
X1066 11847 11928 11931 1 3 NAND2X2 $T=2294160 1380400 0 0 $X=2294158 $Y=1379998
X1067 11927 11615 12040 1 3 NAND2X2 $T=2305380 1299760 0 180 $X=2302080 $Y=1294320
X1068 12043 617 11853 1 3 NAND2X2 $T=2303400 1420720 1 0 $X=2303398 $Y=1415280
X1069 630 12434 12216 1 3 NAND2X2 $T=2366760 1370320 1 0 $X=2366758 $Y=1364880
X1070 12498 12595 12536 1 3 NAND2X2 $T=2389200 1400560 0 0 $X=2389198 $Y=1400158
X1071 641 12957 12928 1 3 NAND2X2 $T=2440020 1340080 1 180 $X=2436720 $Y=1339678
X1072 12999 12908 13064 1 3 NAND2X2 $T=2450580 1330000 0 0 $X=2450578 $Y=1329598
X1073 13277 13272 655 1 3 NAND2X2 $T=2488200 1148560 0 180 $X=2484900 $Y=1143120
X1074 13159 13275 13224 1 3 NAND2X2 $T=2486880 1259440 0 0 $X=2486878 $Y=1259038
X1075 656 13319 13335 1 3 NAND2X2 $T=2496780 1309840 1 0 $X=2496778 $Y=1304400
X1076 13222 13514 13507 1 3 NAND2X2 $T=2514600 1219120 0 180 $X=2511300 $Y=1213680
X1077 664 13561 13348 1 3 NAND2X2 $T=2519220 1269520 1 0 $X=2519218 $Y=1264080
X1078 13701 668 13504 1 3 NAND2X2 $T=2534400 1239280 1 0 $X=2534398 $Y=1233840
X1079 13881 678 13638 1 3 NAND2X2 $T=2552880 1229200 1 0 $X=2552878 $Y=1223760
X1080 677 13929 13424 1 3 NAND2X2 $T=2557500 1209040 1 0 $X=2557498 $Y=1203600
X1081 2893 3 2819 2896 1 2916 AOI21X4 $T=873840 1269520 1 0 $X=873838 $Y=1264080
X1082 2868 3 2941 2977 1 3068 AOI21X4 $T=887700 1198960 0 0 $X=887698 $Y=1198558
X1083 3019 3 3060 3014 1 2978 AOI21X4 $T=903540 1350160 0 180 $X=896940 $Y=1344720
X1084 118 3 3070 3061 1 3023 AOI21X4 $T=908160 1400560 1 180 $X=901560 $Y=1400158
X1085 117 3 3162 3142 1 3113 AOI21X4 $T=926640 1168720 1 180 $X=920040 $Y=1168318
X1086 3371 3 3373 3354 1 3353 AOI21X4 $T=958320 1239280 0 180 $X=951720 $Y=1233840
X1087 3236 3 3358 3378 1 3382 AOI21X4 $T=952380 1309840 0 0 $X=952378 $Y=1309438
X1088 3420 3 3409 3419 1 3297 AOI21X4 $T=968880 1350160 1 180 $X=962280 $Y=1349758
X1089 3708 3 3736 3750 1 3740 AOI21X4 $T=1009800 1319920 0 0 $X=1009798 $Y=1319518
X1090 4051 3 4050 4028 1 3868 AOI21X4 $T=1057320 1400560 1 180 $X=1050720 $Y=1400158
X1091 6309 3 6341 6308 1 6423 AOI21X4 $T=1419660 1239280 1 0 $X=1419658 $Y=1233840
X1092 6481 3 312 6439 1 6506 AOI21X4 $T=1441440 1400560 1 0 $X=1441438 $Y=1395120
X1093 6656 3 6572 6632 1 6672 AOI21X4 $T=1462560 1340080 0 0 $X=1462558 $Y=1339678
X1094 6773 3 6768 6788 1 6946 AOI21X4 $T=1483020 1209040 1 0 $X=1483018 $Y=1203600
X1095 6796 3 6727 6755 1 6855 AOI21X4 $T=1486320 1289680 1 0 $X=1486318 $Y=1284240
X1096 7055 3 6973 7065 1 7073 AOI21X4 $T=1524600 1390480 0 0 $X=1524598 $Y=1390078
X1097 7320 3 7089 7325 1 7329 AOI21X4 $T=1558920 1319920 0 0 $X=1558918 $Y=1319518
X1098 7285 3 7386 7381 1 7522 AOI21X4 $T=1574100 1178800 1 0 $X=1574098 $Y=1173360
X1099 7549 3 7392 7511 1 7520 AOI21X4 $T=1601820 1299760 0 180 $X=1595220 $Y=1294320
X1100 7071 3 7547 7501 1 353 AOI21X4 $T=1604460 1138480 0 0 $X=1604458 $Y=1138078
X1101 7708 3 7658 7686 1 7869 AOI21X4 $T=1624920 1239280 1 0 $X=1624918 $Y=1233840
X1102 7986 3 7959 8008 1 371 AOI21X4 $T=1663200 1168720 1 0 $X=1663198 $Y=1163280
X1103 8894 3 8864 8954 1 8945 AOI21X4 $T=1815000 1350160 1 0 $X=1814998 $Y=1344720
X1104 451 3 9012 9003 1 9069 AOI21X4 $T=1833480 1380400 1 0 $X=1833478 $Y=1374960
X1105 9235 3 9314 9206 1 483 AOI21X4 $T=1876380 1158640 1 0 $X=1876378 $Y=1153200
X1106 9960 3 9920 9959 1 10005 AOI21X4 $T=1980000 1350160 0 0 $X=1979998 $Y=1349758
X1107 10003 3 524 10010 1 10009 AOI21X4 $T=1980660 1319920 1 0 $X=1980658 $Y=1314480
X1108 10076 3 10141 10147 1 10176 AOI21X4 $T=1997820 1279600 0 0 $X=1997818 $Y=1279198
X1109 11849 3 11928 11937 1 11944 AOI21X4 $T=2290200 1390480 1 0 $X=2290198 $Y=1385040
X1110 11964 3 12373 12375 1 12393 AOI21X4 $T=2350920 1360240 0 0 $X=2350918 $Y=1359838
X1111 12247 3 12272 12374 1 12436 AOI21X4 $T=2356200 1269520 1 0 $X=2356198 $Y=1264080
X1112 12565 3 12572 12558 1 634 AOI21X4 $T=2389200 1219120 1 180 $X=2382600 $Y=1218718
X1113 12811 3 12540 12843 1 13156 AOI21X4 $T=2428140 1370320 1 0 $X=2428138 $Y=1364880
X1114 12600 3 12908 12929 1 12902 AOI21X4 $T=2432100 1319920 0 0 $X=2432098 $Y=1319518
X1115 13096 3 13207 13239 1 13244 AOI21X4 $T=2482920 1350160 1 0 $X=2482918 $Y=1344720
X1116 13275 3 13187 13301 1 13240 AOI21X4 $T=2486880 1269520 1 0 $X=2486878 $Y=1264080
X1117 13038 3 13334 13347 1 13458 AOI21X4 $T=2494800 1249360 1 0 $X=2494798 $Y=1243920
X1118 14089 3 13698 14118 1 13941 AOI21X4 $T=2587200 1279600 1 0 $X=2587198 $Y=1274160
X1119 1606 3 1566 1 1600 AND2X2 $T=687060 1239280 1 180 $X=684420 $Y=1238878
X1120 1848 3 1841 1 1633 AND2X2 $T=721380 1340080 1 180 $X=718740 $Y=1339678
X1121 1782 3 1848 1 1749 AND2X2 $T=721380 1360240 0 180 $X=718740 $Y=1354800
X1122 2110 3 2235 1 1993 AND2X2 $T=752400 1299760 0 180 $X=749760 $Y=1294320
X1123 2766 3 2672 1 2817 AND2X2 $T=852720 1209040 1 0 $X=852718 $Y=1203600
X1124 2843 3 2635 1 2789 AND2X2 $T=863940 1178800 1 180 $X=861300 $Y=1178398
X1125 3065 3 3062 1 3069 AND2X2 $T=904200 1390480 1 0 $X=904198 $Y=1385040
X1126 3407 3 134 1 3415 AND2X2 $T=961620 1198960 1 0 $X=961618 $Y=1193520
X1127 3358 3 3437 1 3269 AND2X2 $T=969540 1309840 0 180 $X=966900 $Y=1304400
X1128 3436 3 3445 1 3467 AND2X2 $T=968220 1400560 0 0 $X=968218 $Y=1400158
X1129 130 3 128 1 3464 AND2X2 $T=978120 1219120 0 180 $X=975480 $Y=1213680
X1130 3794 3 3801 1 3805 AND2X2 $T=1021680 1289680 1 0 $X=1021678 $Y=1284240
X1131 212 3 206 1 4538 AND2X2 $T=1145100 1420720 0 0 $X=1145098 $Y=1420318
X1132 187 3 188 1 4947 AND2X2 $T=1206480 1219120 0 180 $X=1203840 $Y=1213680
X1133 259 3 230 1 5374 AND2X2 $T=1254660 1380400 0 0 $X=1254658 $Y=1379998
X1134 6458 3 6433 1 6482 AND2X2 $T=1437480 1289680 1 0 $X=1437478 $Y=1284240
X1135 6440 3 6493 1 313 AND2X2 $T=1445400 1420720 0 0 $X=1445398 $Y=1420318
X1136 6591 3 6278 1 6599 AND2X2 $T=1455960 1188880 0 0 $X=1455958 $Y=1188478
X1137 312 3 6597 1 6637 AND2X2 $T=1461240 1410640 1 0 $X=1461238 $Y=1405200
X1138 6440 3 6676 1 319 AND2X2 $T=1469160 1420720 0 0 $X=1469158 $Y=1420318
X1139 6733 3 6753 1 6802 AND2X2 $T=1482360 1299760 0 0 $X=1482358 $Y=1299358
X1140 6702 3 6792 1 6877 AND2X2 $T=1494240 1168720 0 0 $X=1494238 $Y=1168318
X1141 326 3 325 1 6806 AND2X2 $T=1499520 1420720 1 180 $X=1496880 $Y=1420318
X1142 6798 3 6940 1 6975 AND2X2 $T=1505460 1340080 0 0 $X=1505458 $Y=1339678
X1143 6440 3 6974 1 6821 AND2X2 $T=1512060 1420720 1 180 $X=1509420 $Y=1420318
X1144 332 3 330 1 7066 AND2X2 $T=1521300 1138480 0 0 $X=1521298 $Y=1138078
X1145 7127 3 7027 1 7172 AND2X2 $T=1539780 1249360 1 0 $X=1539778 $Y=1243920
X1146 7285 3 7255 1 7421 AND2X2 $T=1573440 1188880 1 0 $X=1573438 $Y=1183440
X1147 7599 3 7377 1 7675 AND2X2 $T=1620960 1158640 0 0 $X=1620958 $Y=1158238
X1148 8310 3 8309 1 8295 AND2X2 $T=1712700 1148560 0 180 $X=1710060 $Y=1143120
X1149 436 3 432 1 438 AND2X2 $T=1790580 1420720 0 0 $X=1790578 $Y=1420318
X1150 8884 3 8918 1 444 AND2X2 $T=1806420 1400560 1 180 $X=1803780 $Y=1400158
X1151 8922 3 8884 1 450 AND2X2 $T=1814340 1410640 0 180 $X=1811700 $Y=1405200
X1152 440 3 422 1 9065 AND2X2 $T=1822260 1410640 1 0 $X=1822258 $Y=1405200
X1153 436 3 9066 1 9036 AND2X2 $T=1836780 1420720 0 180 $X=1834140 $Y=1415280
X1154 436 3 9070 1 9103 AND2X2 $T=1838100 1410640 1 0 $X=1838098 $Y=1405200
X1155 8884 3 9240 1 9033 AND2X2 $T=1857240 1410640 0 180 $X=1854600 $Y=1405200
X1156 8884 3 9245 1 9122 AND2X2 $T=1861200 1400560 1 180 $X=1858560 $Y=1400158
X1157 9355 3 9381 1 9322 AND2X2 $T=1886280 1380400 0 180 $X=1883640 $Y=1374960
X1158 9533 3 9529 1 9537 AND2X2 $T=1906080 1299760 0 0 $X=1906078 $Y=1299358
X1159 9593 3 9567 1 9631 AND2X2 $T=1921920 1209040 0 0 $X=1921918 $Y=1208638
X1160 9506 3 493 1 9687 AND2X2 $T=1929180 1188880 0 0 $X=1929178 $Y=1188478
X1161 9683 3 435 1 9736 AND2X2 $T=1937100 1209040 1 0 $X=1937098 $Y=1203600
X1162 9855 3 449 1 9739 AND2X2 $T=1955580 1259440 0 180 $X=1952940 $Y=1254000
X1163 10272 3 10270 1 10142 AND2X2 $T=2022240 1299760 0 180 $X=2019600 $Y=1294320
X1164 538 3 10322 1 10384 AND2X2 $T=2065800 1148560 0 180 $X=2063160 $Y=1143120
X1165 10818 3 10820 1 10768 AND2X2 $T=2112660 1400560 1 180 $X=2110020 $Y=1400158
X1166 11821 3 12102 1 12127 AND2X2 $T=2313960 1198960 1 0 $X=2313958 $Y=1193520
X1167 12457 3 12426 1 12293 AND2X2 $T=2367420 1350160 0 180 $X=2364780 $Y=1344720
X1168 12560 3 12286 1 12599 AND2X2 $T=2384580 1239280 0 0 $X=2384578 $Y=1238878
X1169 12746 3 12715 1 12803 AND2X2 $T=2413620 1219120 0 0 $X=2413618 $Y=1218718
X1170 12908 3 12928 1 12629 AND2X2 $T=2435400 1330000 1 180 $X=2432760 $Y=1329598
X1171 13159 3 13090 1 13098 AND2X2 $T=2469720 1269520 0 180 $X=2467080 $Y=1264080
X1172 13207 3 13216 1 13095 AND2X2 $T=2473680 1350160 0 180 $X=2471040 $Y=1344720
X1173 13418 3 13222 1 13427 AND2X2 $T=2502060 1198960 0 0 $X=2502058 $Y=1198558
X1174 13514 3 13504 1 13245 AND2X2 $T=2513940 1229200 1 180 $X=2511300 $Y=1228798
X1175 14035 3 13899 1 13940 AND2X2 $T=2575320 1279600 0 180 $X=2572680 $Y=1274160
X1176 14232 3 14229 1 14078 AND2X2 $T=2604360 1229200 1 180 $X=2601720 $Y=1228798
X1177 53 1 2947 3 2946 NAND2X4 $T=889020 1279600 0 0 $X=889018 $Y=1279198
X1178 7653 1 6950 3 7650 NAND2X4 $T=1615020 1259440 1 180 $X=1610400 $Y=1259038
X1179 7600 1 366 3 7987 NAND2X4 $T=1665840 1188880 0 0 $X=1665838 $Y=1188478
X1180 476 1 475 3 9101 NAND2X4 $T=1866480 1168720 1 180 $X=1861860 $Y=1168318
X1181 9350 1 9317 3 9235 NAND2X4 $T=1879680 1370320 1 180 $X=1875060 $Y=1369918
X1182 9868 1 9848 3 9536 NAND2X4 $T=1952940 1309840 0 180 $X=1948320 $Y=1304400
X1183 515 1 513 3 9668 NAND2X4 $T=1955580 1319920 1 180 $X=1950960 $Y=1319518
X1184 9868 1 9880 3 9872 NAND2X4 $T=1957560 1269520 0 0 $X=1957558 $Y=1269118
X1185 9903 1 9960 3 9985 NAND2X4 $T=1980000 1360240 1 0 $X=1979998 $Y=1354800
X1186 10143 1 10076 3 10174 NAND2X4 $T=2008380 1279600 0 0 $X=2008378 $Y=1279198
X1187 11554 1 11549 3 6948 NAND2X4 $T=2235420 1390480 1 180 $X=2230800 $Y=1390078
X1188 13188 1 650 3 13090 NAND2X4 $T=2473680 1279600 0 0 $X=2473678 $Y=1279198
X1189 62 58 1 3 1509 OR2X2 $T=665940 1249360 1 0 $X=665938 $Y=1243920
X1190 55 1748 1 3 1814 OR2X2 $T=708180 1249360 0 0 $X=708178 $Y=1248958
X1191 76 1842 1 3 1787 OR2X2 $T=720060 1430800 0 180 $X=717420 $Y=1425360
X1192 1918 1842 1 3 1849 OR2X2 $T=727980 1430800 0 180 $X=725340 $Y=1425360
X1193 1806 1915 1 3 1847 OR2X2 $T=729300 1269520 0 180 $X=726660 $Y=1264080
X1194 1898 1956 1 3 1943 OR2X2 $T=736560 1360240 1 180 $X=733920 $Y=1359838
X1195 1923 82 1 3 1985 OR2X2 $T=736560 1178800 1 0 $X=736558 $Y=1173360
X1196 2251 2214 1 3 2138 OR2X2 $T=770880 1178800 0 180 $X=768240 $Y=1173360
X1197 2281 2321 1 3 2237 OR2X2 $T=786060 1279600 0 180 $X=783420 $Y=1274160
X1198 2370 2374 1 3 2241 OR2X2 $T=793320 1239280 0 180 $X=790680 $Y=1233840
X1199 2330 2341 1 3 2305 OR2X2 $T=794640 1219120 0 180 $X=792000 $Y=1213680
X1200 92 93 1 3 94 OR2X2 $T=793320 1148560 1 0 $X=793318 $Y=1143120
X1201 87 99 1 3 2269 OR2X2 $T=823020 1178800 1 180 $X=820380 $Y=1178398
X1202 95 101 1 3 2490 OR2X2 $T=823020 1420720 0 180 $X=820380 $Y=1415280
X1203 3192 3089 1 3 3171 OR2X2 $T=928620 1390480 1 180 $X=925980 $Y=1390078
X1204 125 3266 1 3 3162 OR2X2 $T=944460 1178800 0 180 $X=941820 $Y=1173360
X1205 3349 126 1 3 3137 OR2X2 $T=945780 1158640 0 180 $X=943140 $Y=1153200
X1206 3534 137 1 3 3409 OR2X2 $T=969540 1360240 0 180 $X=966900 $Y=1354800
X1207 3505 3550 1 3 3408 OR2X2 $T=989340 1410640 1 180 $X=986700 $Y=1410238
X1208 158 3731 1 3 3713 OR2X2 $T=1011120 1420720 0 180 $X=1008480 $Y=1415280
X1209 3951 4021 1 3 3856 OR2X2 $T=1051380 1360240 1 180 $X=1048740 $Y=1359838
X1210 4093 4089 1 3 3857 OR2X2 $T=1063920 1370320 1 180 $X=1061280 $Y=1369918
X1211 4186 4215 1 3 173 OR2X2 $T=1087020 1420720 0 180 $X=1084380 $Y=1415280
X1212 192 198 1 3 4306 OR2X2 $T=1112100 1340080 0 180 $X=1109460 $Y=1334640
X1213 188 5108 1 3 5266 OR2X2 $T=1230900 1249360 0 0 $X=1230898 $Y=1248958
X1214 101 5465 1 3 5486 OR2X2 $T=1275780 1330000 0 0 $X=1275778 $Y=1329598
X1215 5521 265 1 3 5465 OR2X2 $T=1279740 1350160 1 180 $X=1277100 $Y=1349758
X1216 97 5555 1 3 5571 OR2X2 $T=1290960 1319920 0 0 $X=1290958 $Y=1319518
X1217 104 5576 1 3 5654 OR2X2 $T=1293600 1249360 1 0 $X=1293598 $Y=1243920
X1218 110 5571 1 3 5585 OR2X2 $T=1293600 1299760 0 0 $X=1293598 $Y=1299358
X1219 235 5585 1 3 5576 OR2X2 $T=1296900 1279600 1 180 $X=1294260 $Y=1279198
X1220 264 5587 1 3 5521 OR2X2 $T=1296900 1360240 0 180 $X=1294260 $Y=1354800
X1221 108 5586 1 3 286 OR2X2 $T=1333200 1209040 0 0 $X=1333198 $Y=1208638
X1222 288 284 1 3 5922 OR2X2 $T=1341120 1360240 1 0 $X=1341118 $Y=1354800
X1223 6000 5997 1 3 6088 OR2X2 $T=1370160 1330000 1 0 $X=1370158 $Y=1324560
X1224 6039 6068 1 3 6095 OR2X2 $T=1377420 1319920 1 0 $X=1377418 $Y=1314480
X1225 6277 6165 1 3 6422 OR2X2 $T=1413060 1198960 1 0 $X=1413058 $Y=1193520
X1226 6335 6160 1 3 6405 OR2X2 $T=1422960 1168720 0 0 $X=1422958 $Y=1168318
X1227 6378 5711 1 3 6458 OR2X2 $T=1426260 1279600 0 0 $X=1426258 $Y=1279198
X1228 6637 6628 1 3 6675 OR2X2 $T=1463880 1410640 1 0 $X=1463878 $Y=1405200
X1229 3093 320 1 3 6733 OR2X2 $T=1475760 1299760 1 0 $X=1475758 $Y=1294320
X1230 6695 6693 1 3 6737 OR2X2 $T=1477080 1148560 0 0 $X=1477078 $Y=1148158
X1231 3352 322 1 3 6798 OR2X2 $T=1487640 1340080 0 0 $X=1487638 $Y=1339678
X1232 6948 6941 1 3 6920 OR2X2 $T=1510740 1390480 0 180 $X=1508100 $Y=1385040
X1233 7005 3355 1 3 7127 OR2X2 $T=1519320 1259440 0 180 $X=1516680 $Y=1254000
X1234 7138 337 1 3 7282 OR2X2 $T=1555620 1269520 0 0 $X=1555618 $Y=1269118
X1235 337 335 1 3 7283 OR2X2 $T=1555620 1279600 1 0 $X=1555618 $Y=1274160
X1236 7282 7349 1 3 7328 OR2X2 $T=1570800 1249360 1 180 $X=1568160 $Y=1248958
X1237 7283 338 1 3 7379 OR2X2 $T=1570140 1279600 1 0 $X=1570138 $Y=1274160
X1238 7384 7282 1 3 7358 OR2X2 $T=1574100 1239280 1 180 $X=1571460 $Y=1238878
X1239 7177 7502 1 3 7604 OR2X2 $T=1592580 1319920 0 0 $X=1592578 $Y=1319518
X1240 7801 356 1 3 7790 OR2X2 $T=1640100 1410640 1 180 $X=1637460 $Y=1410238
X1241 6671 8168 1 3 8245 OR2X2 $T=1695540 1309840 1 0 $X=1695538 $Y=1304400
X1242 8166 8172 1 3 8175 OR2X2 $T=1696200 1209040 1 0 $X=1696198 $Y=1203600
X1243 8188 8240 1 3 8249 OR2X2 $T=1698840 1209040 1 0 $X=1698838 $Y=1203600
X1244 6568 8574 1 3 8496 OR2X2 $T=1754280 1289680 1 180 $X=1751640 $Y=1289278
X1245 7352 8656 1 3 8731 OR2X2 $T=1775400 1188880 0 0 $X=1775398 $Y=1188478
X1246 7010 8627 1 3 8653 OR2X2 $T=1775400 1209040 0 0 $X=1775398 $Y=1208638
X1247 6825 8863 1 3 8749 OR2X2 $T=1802460 1239280 0 0 $X=1802458 $Y=1238878
X1248 491 492 1 3 9355 OR2X2 $T=1904760 1370320 1 180 $X=1902120 $Y=1369918
X1249 8780 9764 1 3 9757 OR2X2 $T=1944360 1239280 1 180 $X=1941720 $Y=1238878
X1250 9791 9780 1 3 9773 OR2X2 $T=1947000 1239280 1 180 $X=1944360 $Y=1238878
X1251 521 511 1 3 9814 OR2X2 $T=1952940 1350160 1 180 $X=1950300 $Y=1349758
X1252 508 9696 1 3 9851 OR2X2 $T=1950960 1410640 1 0 $X=1950958 $Y=1405200
X1253 9812 9791 1 3 9867 OR2X2 $T=1952280 1229200 0 0 $X=1952278 $Y=1228798
X1254 519 9895 1 3 9900 OR2X2 $T=1960860 1410640 0 0 $X=1960858 $Y=1410238
X1255 520 9722 1 3 9895 OR2X2 $T=1960860 1420720 1 0 $X=1960858 $Y=1415280
X1256 8780 9929 1 3 9871 OR2X2 $T=1971420 1229200 1 180 $X=1968780 $Y=1228798
X1257 523 10177 1 3 10171 OR2X2 $T=2010360 1400560 0 180 $X=2007720 $Y=1395120
X1258 10264 10174 1 3 10203 OR2X2 $T=2018280 1309840 0 180 $X=2015640 $Y=1304400
X1259 518 520 1 3 10421 OR2X2 $T=2038080 1390480 0 0 $X=2038078 $Y=1390078
X1260 548 10387 1 3 10268 OR2X2 $T=2046000 1420720 1 180 $X=2043360 $Y=1420318
X1261 538 10322 1 3 547 OR2X2 $T=2055900 1138480 1 180 $X=2053260 $Y=1138078
X1262 550 552 1 3 10387 OR2X2 $T=2057880 1420720 0 0 $X=2057878 $Y=1420318
X1263 10432 10496 1 3 541 OR2X2 $T=2060520 1148560 1 180 $X=2057880 $Y=1148158
X1264 10480 10476 1 3 10501 OR2X2 $T=2065800 1259440 1 0 $X=2065798 $Y=1254000
X1265 555 549 1 3 10623 OR2X2 $T=2082300 1400560 1 0 $X=2082298 $Y=1395120
X1266 579 10784 1 3 10818 OR2X2 $T=2107380 1410640 0 0 $X=2107378 $Y=1410238
X1267 10860 10820 1 3 10821 OR2X2 $T=2116620 1390480 0 180 $X=2113980 $Y=1385040
X1268 10889 10893 1 3 10890 OR2X2 $T=2128500 1400560 1 180 $X=2125860 $Y=1400158
X1269 570 10172 1 3 11030 OR2X2 $T=2142360 1380400 0 0 $X=2142358 $Y=1379998
X1270 11071 592 1 3 11128 OR2X2 $T=2159520 1420720 0 0 $X=2159518 $Y=1420318
X1271 9851 604 1 3 605 OR2X2 $T=2199780 1198960 0 0 $X=2199778 $Y=1198558
X1272 11908 12212 1 3 12372 OR2X2 $T=2350260 1168720 1 0 $X=2350258 $Y=1163280
X1273 12477 12326 1 3 12498 OR2X2 $T=2374020 1400560 1 0 $X=2374018 $Y=1395120
X1274 641 12957 1 3 12908 OR2X2 $T=2440020 1330000 0 0 $X=2440018 $Y=1329598
X1275 13218 12939 1 3 13207 OR2X2 $T=2485560 1350160 0 0 $X=2485558 $Y=1349758
X1276 13287 13279 1 3 13273 OR2X2 $T=2489520 1188880 1 180 $X=2486880 $Y=1188478
X1277 651 13305 1 3 13277 OR2X2 $T=2495460 1158640 0 180 $X=2492820 $Y=1153200
X1278 13461 12844 1 3 13501 OR2X2 $T=2507340 1330000 0 0 $X=2507338 $Y=1329598
X1279 13785 13774 1 3 13457 OR2X2 $T=2545620 1178800 1 180 $X=2542980 $Y=1178398
X1280 672 670 1 3 13816 OR2X2 $T=2549580 1430800 0 180 $X=2546940 $Y=1425360
X1281 13882 12870 1 3 13814 OR2X2 $T=2554860 1309840 0 180 $X=2552220 $Y=1304400
X1282 13987 13971 1 3 13913 OR2X2 $T=2570040 1370320 0 180 $X=2567400 $Y=1364880
X1283 675 688 1 3 13900 OR2X2 $T=2580600 1380400 1 180 $X=2577960 $Y=1379998
X1284 693 692 1 3 14139 OR2X2 $T=2599080 1410640 1 180 $X=2596440 $Y=1410238
X1285 1782 1 3 1750 1658 NAND2XL $T=702240 1370320 1 180 $X=700260 $Y=1369918
X1286 1749 1 3 1750 1754 NAND2XL $T=702900 1360240 1 0 $X=702898 $Y=1354800
X1287 1917 1 3 1815 1701 NAND2XL $T=723360 1420720 0 180 $X=721380 $Y=1415280
X1288 82 1 3 1923 1927 NAND2XL $T=729300 1178800 1 0 $X=729298 $Y=1173360
X1289 2177 1 3 2110 2172 NAND2XL $T=764940 1279600 1 180 $X=762960 $Y=1279198
X1290 2271 1 3 2212 2251 NAND2XL $T=776820 1188880 0 180 $X=774840 $Y=1183440
X1291 2342 1 3 2336 1841 NAND2XL $T=787380 1340080 1 180 $X=785400 $Y=1339678
X1292 2316 1 3 2212 2368 NAND2XL $T=789360 1188880 0 0 $X=789358 $Y=1188478
X1293 3435 1 3 3409 3406 NAND2XL $T=962940 1360240 0 180 $X=960960 $Y=1354800
X1294 169 1 3 3674 3589 NAND2XL $T=1025640 1148560 1 180 $X=1023660 $Y=1148158
X1295 166 1 3 165 3731 NAND2XL $T=1026960 1420720 0 180 $X=1024980 $Y=1415280
X1296 4086 1 3 4060 4061 NAND2XL $T=1065900 1188880 0 180 $X=1063920 $Y=1183440
X1297 4209 1 3 4149 4177 NAND2XL $T=1081740 1269520 1 180 $X=1079760 $Y=1269118
X1298 187 1 3 191 4262 NAND2XL $T=1098900 1420720 1 180 $X=1096920 $Y=1420318
X1299 191 1 3 189 4267 NAND2XL $T=1102860 1410640 1 180 $X=1100880 $Y=1410238
X1300 187 1 3 189 4265 NAND2XL $T=1115400 1420720 0 180 $X=1113420 $Y=1415280
X1301 4367 1 3 4460 4439 NAND2XL $T=1131240 1319920 1 180 $X=1129260 $Y=1319518
X1302 186 1 3 210 5757 NAND2XL $T=1319340 1330000 1 0 $X=1319338 $Y=1324560
X1303 6763 1 3 6759 6820 NAND2XL $T=1487640 1330000 0 0 $X=1487638 $Y=1329598
X1304 6944 1 3 6920 6880 NAND2XL $T=1505460 1390480 1 180 $X=1503480 $Y=1390078
X1305 7074 1 3 7103 7160 NAND2XL $T=1539780 1360240 1 0 $X=1539778 $Y=1354800
X1306 7056 1 3 7055 7262 NAND2XL $T=1550340 1400560 0 0 $X=1550338 $Y=1400158
X1307 7214 1 3 7292 7326 NAND2XL $T=1566180 1370320 0 0 $X=1566178 $Y=1369918
X1308 7471 1 3 7392 7603 NAND2XL $T=1592580 1309840 1 0 $X=1592578 $Y=1304400
X1309 7543 1 3 7604 7647 NAND2XL $T=1605120 1309840 0 0 $X=1605118 $Y=1309438
X1310 7837 1 3 7765 7826 NAND2XL $T=1644060 1219120 0 180 $X=1642080 $Y=1213680
X1311 7797 1 3 7764 7918 NAND2XL $T=1647360 1239280 1 0 $X=1647358 $Y=1233840
X1312 8149 1 3 8145 8164 NAND2XL $T=1693560 1239280 0 180 $X=1691580 $Y=1233840
X1313 8100 1 3 8154 381 NAND2XL $T=1692900 1370320 0 0 $X=1692898 $Y=1369918
X1314 8173 1 3 6666 8266 NAND2XL $T=1696860 1340080 0 0 $X=1696858 $Y=1339678
X1315 8243 1 3 8245 8267 NAND2XL $T=1699500 1309840 0 0 $X=1699498 $Y=1309438
X1316 8242 1 3 387 8241 NAND2XL $T=1712040 1239280 0 180 $X=1710060 $Y=1233840
X1317 8149 1 3 8368 8401 NAND2XL $T=1727880 1168720 0 0 $X=1727878 $Y=1168318
X1318 8373 1 3 387 8452 NAND2XL $T=1731180 1168720 0 0 $X=1731178 $Y=1168318
X1319 8477 1 3 8496 8495 NAND2XL $T=1747680 1289680 0 180 $X=1745700 $Y=1284240
X1320 8633 1 3 8653 8707 NAND2XL $T=1767480 1219120 1 0 $X=1767478 $Y=1213680
X1321 8658 1 3 8731 8759 NAND2XL $T=1783320 1188880 0 0 $X=1783318 $Y=1188478
X1322 8729 1 3 8749 8754 NAND2XL $T=1787280 1249360 1 0 $X=1787278 $Y=1243920
X1323 8861 1 3 8807 8858 NAND2XL $T=1799820 1370320 0 180 $X=1797840 $Y=1364880
X1324 8892 1 3 8886 8890 NAND2XL $T=1809060 1188880 0 180 $X=1807080 $Y=1183440
X1325 8916 1 3 8894 8889 NAND2XL $T=1809060 1350160 1 180 $X=1807080 $Y=1349758
X1326 9383 1 3 9381 9325 NAND2XL $T=1890240 1400560 1 180 $X=1888260 $Y=1400158
X1327 9438 1 3 9355 9360 NAND2XL $T=1896180 1380400 0 180 $X=1894200 $Y=1374960
X1328 9665 1 3 9632 9628 NAND2XL $T=1923900 1340080 1 180 $X=1921920 $Y=1339678
X1329 9668 1 3 9689 9713 NAND2XL $T=1935120 1319920 0 0 $X=1935118 $Y=1319518
X1330 10170 1 3 10076 10052 NAND2XL $T=1999800 1269520 1 180 $X=1997820 $Y=1269118
X1331 10051 1 3 10143 10011 NAND2XL $T=2000460 1269520 1 0 $X=2000458 $Y=1264080
X1332 10396 1 3 541 10274 NAND2XL $T=2042700 1148560 1 180 $X=2040720 $Y=1148158
X1333 556 1 3 10497 10357 NAND2XL $T=2066460 1360240 0 180 $X=2064480 $Y=1354800
X1334 11579 1 3 11734 11549 NAND2XL $T=2251920 1390480 1 180 $X=2249940 $Y=1390078
X1335 12041 1 3 11928 11874 NAND2XL $T=2303400 1390480 0 180 $X=2301420 $Y=1385040
X1336 621 1 3 11965 12276 NAND2XL $T=2323200 1138480 0 0 $X=2323198 $Y=1138078
X1337 12286 1 3 12496 12500 NAND2XL $T=2374680 1239280 0 0 $X=2374678 $Y=1238878
X1338 12325 1 3 12372 12564 NAND2XL $T=2382600 1168720 0 0 $X=2382598 $Y=1168318
X1339 12292 1 3 12622 12743 NAND2XL $T=2403720 1198960 0 0 $X=2403718 $Y=1198558
X1340 609 1 3 12042 12818 NAND2XL $T=2409660 1168720 1 0 $X=2409658 $Y=1163280
X1341 12835 1 3 638 12903 NAND2XL $T=2431440 1158640 1 0 $X=2431438 $Y=1153200
X1342 647 1 3 13092 12993 NAND2XL $T=2457840 1400560 0 180 $X=2455860 $Y=1395120
X1343 13092 1 3 13088 13087 NAND2XL $T=2458500 1420720 1 180 $X=2456520 $Y=1420318
X1344 13335 1 3 13275 13000 NAND2XL $T=2494140 1279600 0 180 $X=2492160 $Y=1274160
X1345 13501 1 3 13500 13270 NAND2XL $T=2512620 1340080 0 180 $X=2510640 $Y=1334640
X1346 13552 1 3 13088 13562 NAND2XL $T=2518560 1420720 1 0 $X=2518558 $Y=1415280
X1347 13651 1 3 13684 13696 NAND2XL $T=2532420 1400560 0 0 $X=2532418 $Y=1400158
X1348 13122 1 3 13769 13790 NAND2XL $T=2542980 1168720 1 0 $X=2542978 $Y=1163280
X1349 679 1 3 13985 13949 NAND2XL $T=2570700 1148560 1 0 $X=2570698 $Y=1143120
X1350 682 1 3 683 13946 NAND2XL $T=2572680 1410640 1 180 $X=2570700 $Y=1410238
X1351 14143 1 3 14090 13987 NAND2XL $T=2588520 1370320 1 180 $X=2586540 $Y=1369918
X1352 696 1 3 14090 14312 NAND2XL $T=2611620 1400560 0 0 $X=2611618 $Y=1400158
X1353 14311 1 3 14090 14280 NAND2XL $T=2616900 1370320 1 180 $X=2614920 $Y=1369918
X1354 57 55 1 3 INVX4 $T=663300 1319920 0 180 $X=660660 $Y=1314480
X1355 1508 62 1 3 INVX4 $T=667260 1309840 0 0 $X=667258 $Y=1309438
X1356 72 76 1 3 INVX4 $T=718740 1400560 1 180 $X=716100 $Y=1400158
X1357 2893 2954 1 3 INVX4 $T=891000 1259440 1 180 $X=888360 $Y=1259038
X1358 3297 3236 1 3 INVX4 $T=948420 1309840 0 180 $X=945780 $Y=1304400
X1359 3740 3732 1 3 INVX4 $T=1011780 1279600 0 180 $X=1009140 $Y=1274160
X1360 3868 3816 1 3 INVX4 $T=1032240 1400560 0 180 $X=1029600 $Y=1395120
X1361 4451 189 1 3 INVX4 $T=1127280 1420720 0 0 $X=1127278 $Y=1420318
X1362 189 204 1 3 INVX4 $T=1143120 1168720 1 0 $X=1143118 $Y=1163280
X1363 177 214 1 3 INVX4 $T=1148400 1188880 0 180 $X=1145760 $Y=1183440
X1364 196 199 1 3 INVX4 $T=1173480 1269520 1 0 $X=1173478 $Y=1264080
X1365 187 182 1 3 INVX4 $T=1178100 1239280 0 180 $X=1175460 $Y=1233840
X1366 191 210 1 3 INVX4 $T=1226280 1330000 0 0 $X=1226278 $Y=1329598
X1367 188 186 1 3 INVX4 $T=1249380 1330000 0 180 $X=1246740 $Y=1324560
X1368 6672 6972 1 3 INVX4 $T=1502820 1330000 1 0 $X=1502818 $Y=1324560
X1369 6855 7179 1 3 INVX4 $T=1550340 1239280 0 0 $X=1550338 $Y=1238878
X1370 7178 7285 1 3 INVX4 $T=1558260 1178800 1 0 $X=1558258 $Y=1173360
X1371 7790 7527 1 3 INVX4 $T=1637460 1400560 0 0 $X=1637458 $Y=1400158
X1372 7959 7956 1 3 INVX4 $T=1659900 1209040 0 180 $X=1657260 $Y=1203600
X1373 8780 493 1 3 INVX4 $T=1911360 1289680 0 180 $X=1908720 $Y=1284240
X1374 9986 9960 1 3 INVX4 $T=1979340 1360240 1 180 $X=1976700 $Y=1359838
X1375 10205 551 1 3 INVX4 $T=2058540 1299760 0 180 $X=2055900 $Y=1294320
X1376 562 10529 1 3 INVX4 $T=2122560 1299760 1 0 $X=2122558 $Y=1294320
X1377 10520 567 1 3 INVX4 $T=2148960 1259440 0 0 $X=2148958 $Y=1259038
X1378 10302 570 1 3 INVX4 $T=2180640 1168720 1 180 $X=2178000 $Y=1168318
X1379 11284 11451 1 3 INVX4 $T=2216940 1420720 0 0 $X=2216938 $Y=1420318
X1380 620 618 1 3 INVX4 $T=2320560 1430800 0 180 $X=2317920 $Y=1425360
X1381 11707 12192 1 3 INVX4 $T=2337720 1309840 1 0 $X=2337718 $Y=1304400
X1382 12393 12600 1 3 INVX4 $T=2403060 1319920 0 0 $X=2403058 $Y=1319518
X1383 13038 13094 1 3 INVX4 $T=2463120 1249360 1 180 $X=2460480 $Y=1248958
X1384 13090 13187 1 3 INVX4 $T=2473680 1269520 1 0 $X=2473678 $Y=1264080
X1385 13306 13275 1 3 INVX4 $T=2494140 1289680 0 180 $X=2491500 $Y=1284240
X1386 57 1567 3 1569 1700 1 AOI21X1 $T=677160 1299760 0 0 $X=677158 $Y=1299358
X1387 1744 1597 3 1577 1572 1 AOI21X1 $T=681780 1269520 0 180 $X=679140 $Y=1264080
X1388 1606 1664 3 1656 1629 1 AOI21X1 $T=693660 1249360 0 0 $X=693658 $Y=1248958
X1389 66 1779 3 1780 1773 1 AOI21X1 $T=706860 1239280 1 0 $X=706858 $Y=1233840
X1390 77 1815 3 1817 1821 1 AOI21X1 $T=713460 1420720 1 0 $X=713458 $Y=1415280
X1391 2012 77 3 2018 1916 1 AOI21X1 $T=743160 1410640 1 0 $X=743158 $Y=1405200
X1392 1752 2108 3 2111 1958 1 AOI21X1 $T=751080 1350160 0 0 $X=751078 $Y=1349758
X1393 2241 2270 3 2279 2278 1 AOI21X1 $T=777480 1219120 0 0 $X=777478 $Y=1218718
X1394 3236 3248 3 3252 3264 1 AOI21X1 $T=940500 1309840 1 0 $X=940498 $Y=1304400
X1395 150 3674 3 3734 3739 1 AOI21X1 $T=1009800 1148560 0 0 $X=1009798 $Y=1148158
X1396 3857 3816 3 3861 3864 1 AOI21X1 $T=1030920 1370320 0 0 $X=1030918 $Y=1369918
X1397 173 172 3 4126 4091 1 AOI21X1 $T=1071840 1420720 1 180 $X=1069200 $Y=1420318
X1398 166 216 3 4614 4507 1 AOI21X1 $T=1150380 1420720 1 0 $X=1150378 $Y=1415280
X1399 4988 4989 3 4991 4987 1 AOI21X1 $T=1208460 1360240 1 0 $X=1208458 $Y=1354800
X1400 5032 4986 3 4957 5023 1 AOI21X1 $T=1215720 1148560 0 180 $X=1213080 $Y=1143120
X1401 245 224 3 5071 4988 1 AOI21X1 $T=1218360 1350160 1 0 $X=1218358 $Y=1344720
X1402 191 247 3 188 5109 1 AOI21X1 $T=1222980 1299760 1 0 $X=1222978 $Y=1294320
X1403 198 247 3 4778 253 1 AOI21X1 $T=1238160 1138480 1 180 $X=1235520 $Y=1138078
X1404 247 260 3 5374 5260 1 AOI21X1 $T=1262580 1390480 1 180 $X=1259940 $Y=1390078
X1405 6260 6095 3 6254 6255 1 AOI21X1 $T=1404480 1319920 0 180 $X=1401840 $Y=1314480
X1406 6920 6878 3 6973 7037 1 AOI21X1 $T=1510740 1400560 0 0 $X=1510738 $Y=1400158
X1407 7604 7622 3 7549 7646 1 AOI21X1 $T=1607760 1309840 1 0 $X=1607758 $Y=1304400
X1408 7764 7876 3 7875 7933 1 AOI21X1 $T=1649340 1229200 1 0 $X=1649338 $Y=1223760
X1409 380 8154 3 8147 8150 1 AOI21X1 $T=1695540 1370320 0 180 $X=1692900 $Y=1364880
X1410 382 368 3 383 8246 1 AOI21X1 $T=1698180 1390480 0 0 $X=1698178 $Y=1390078
X1411 8363 8496 3 8488 8491 1 AOI21X1 $T=1747020 1289680 1 180 $X=1744380 $Y=1289278
X1412 8653 8704 3 8682 8752 1 AOI21X1 $T=1782000 1219120 1 0 $X=1781998 $Y=1213680
X1413 8784 8764 3 8792 8782 1 AOI21X1 $T=1793880 1158640 1 0 $X=1793878 $Y=1153200
X1414 9353 9355 3 9359 9350 1 AOI21X1 $T=1883640 1370320 0 0 $X=1883638 $Y=1369918
X1415 9814 9924 3 9920 9899 1 AOI21X1 $T=1970100 1340080 1 180 $X=1967460 $Y=1339678
X1416 541 10275 3 10294 10265 1 AOI21X1 $T=2028840 1148560 1 180 $X=2026200 $Y=1148158
X1417 10392 10629 3 10632 10527 1 AOI21X1 $T=2084940 1319920 1 0 $X=2084938 $Y=1314480
X1418 10863 584 3 10868 10894 1 AOI21X1 $T=2120580 1420720 1 0 $X=2120578 $Y=1415280
X1419 600 11128 3 11180 11179 1 AOI21X1 $T=2178000 1420720 1 180 $X=2175360 $Y=1420318
X1420 11092 11276 3 11279 11284 1 AOI21X1 $T=2191860 1420720 1 0 $X=2191858 $Y=1415280
X1421 12467 12395 3 12433 12431 1 AOI21X1 $T=2367420 1209040 1 180 $X=2364780 $Y=1208638
X1422 12372 12465 3 12462 12460 1 AOI21X1 $T=2370060 1178800 1 180 $X=2367420 $Y=1178398
X1423 12492 12598 3 12395 12721 1 AOI21X1 $T=2403060 1239280 1 0 $X=2403058 $Y=1233840
X1424 12807 12598 3 12773 12778 1 AOI21X1 $T=2416260 1229200 1 180 $X=2413620 $Y=1228798
X1425 13501 13239 3 13509 13502 1 AOI21X1 $T=2511960 1340080 0 0 $X=2511958 $Y=1339678
X1426 13899 13942 3 13939 13930 1 AOI21X1 $T=2566080 1269520 1 180 $X=2563440 $Y=1269118
X1427 679 13950 3 13938 13945 1 AOI21X1 $T=2567400 1148560 1 180 $X=2564760 $Y=1148158
X1428 14143 14010 3 14161 13972 1 AOI21X1 $T=2600400 1370320 1 180 $X=2597760 $Y=1369918
X1429 2842 2689 1 2672 3 2767 OAI21X2 $T=865260 1209040 0 180 $X=859980 $Y=1203600
X1430 2946 2870 1 2937 3 2896 OAI21X2 $T=887040 1269520 1 0 $X=887038 $Y=1264080
X1431 3022 2942 1 2984 3 3014 OAI21X2 $T=898920 1340080 1 0 $X=898918 $Y=1334640
X1432 3707 3695 1 3698 3 3697 OAI21X2 $T=1009140 1249360 0 180 $X=1003860 $Y=1243920
X1433 6753 6699 1 6732 3 6755 OAI21X2 $T=1482360 1289680 0 180 $X=1477080 $Y=1284240
X1434 6575 6664 1 6735 3 6788 OAI21X2 $T=1485000 1209040 1 180 $X=1479720 $Y=1208638
X1435 6635 6769 1 6575 3 6838 OAI21X2 $T=1490280 1229200 0 180 $X=1485000 $Y=1223760
X1436 7324 7278 1 7286 3 7325 OAI21X2 $T=1562880 1330000 1 180 $X=1557600 $Y=1329598
X1437 7542 7632 1 7522 3 7624 OAI21X2 $T=1610400 1178800 0 180 $X=1605120 $Y=1173360
X1438 7987 7932 1 7981 3 8008 OAI21X2 $T=1667820 1178800 1 180 $X=1662540 $Y=1178398
X1439 8491 8590 1 8622 3 8755 OAI21X2 $T=1767480 1279600 0 180 $X=1762200 $Y=1274160
X1440 9101 9208 1 9190 3 9206 OAI21X2 $T=1858560 1158640 0 180 $X=1853280 $Y=1153200
X1441 9703 9894 1 9899 3 9947 OAI21X2 $T=1960860 1330000 0 0 $X=1960858 $Y=1329598
X1442 10009 10036 1 10051 3 10037 OAI21X2 $T=1989900 1269520 1 0 $X=1989898 $Y=1264080
X1443 10264 10176 1 10272 3 10261 OAI21X2 $T=2020920 1309840 1 0 $X=2020918 $Y=1304400
X1444 12286 12396 1 12279 3 12395 OAI21X2 $T=2358180 1229200 1 180 $X=2352900 $Y=1228798
X1445 12399 12216 1 12426 3 12375 OAI21X2 $T=2358180 1350160 0 0 $X=2358178 $Y=1349758
X1446 12522 12436 1 12431 3 12558 OAI21X2 $T=2379300 1229200 0 180 $X=2374020 $Y=1223760
X1447 12505 12192 1 12273 3 12528 OAI21X2 $T=2375340 1279600 0 0 $X=2375338 $Y=1279198
X1448 12717 12632 1 12725 3 12724 OAI21X2 $T=2400420 1370320 1 0 $X=2400418 $Y=1364880
X1449 12725 12777 1 12819 3 12843 OAI21X2 $T=2423520 1370320 0 180 $X=2418240 $Y=1364880
X1450 13224 13094 1 13240 3 13241 OAI21X2 $T=2478960 1249360 0 0 $X=2478958 $Y=1248958
X1451 13515 13156 1 13502 3 13512 OAI21X2 $T=2516580 1360240 0 180 $X=2511300 $Y=1354800
X1452 13504 13645 1 13638 3 13339 OAI21X2 $T=2533080 1219120 0 0 $X=2533078 $Y=1218718
X1453 1701 1693 65 1 3 XNOR2X4 $T=700920 1430800 0 180 $X=689700 $Y=1425360
X1454 112 113 2820 1 3 XNOR2X4 $T=848760 1138480 0 0 $X=848758 $Y=1138078
X1455 3008 3021 3355 1 3 XNOR2X4 $T=897600 1249360 0 0 $X=897598 $Y=1248958
X1456 2817 3068 3246 1 3 XNOR2X4 $T=904200 1209040 1 0 $X=904198 $Y=1203600
X1457 3161 3171 3350 1 3 XNOR2X4 $T=924660 1380400 0 0 $X=924658 $Y=1379998
X1458 2979 3158 3359 1 3 XNOR2X4 $T=932580 1330000 0 0 $X=932578 $Y=1329598
X1459 3405 3382 2939 1 3 XNOR2X4 $T=962280 1319920 1 180 $X=951060 $Y=1319518
X1460 6795 6826 6950 1 3 XNOR2X4 $T=1489620 1269520 0 0 $X=1489618 $Y=1269118
X1461 506 9696 522 1 3 XNOR2X4 $T=1945020 1400560 1 0 $X=1945018 $Y=1395120
X1462 10052 10037 9880 1 3 XNOR2X4 $T=1994520 1269520 1 180 $X=1983300 $Y=1269118
X1463 517 10171 10205 1 3 XNOR2X4 $T=2002440 1410640 1 0 $X=2002438 $Y=1405200
X1464 10235 10231 9848 1 3 XNOR2X4 $T=2018940 1330000 0 180 $X=2007720 $Y=1324560
X1465 11705 11582 613 1 3 XNOR2X4 $T=2250600 1360240 0 0 $X=2250598 $Y=1359838
X1466 12401 12425 12435 1 3 XNOR2X4 $T=2359500 1309840 1 0 $X=2359498 $Y=1304400
X1467 12501 12528 12569 1 3 XNOR2X4 $T=2376000 1289680 1 0 $X=2375998 $Y=1284240
X1468 13000 12992 7597 1 3 XNOR2X4 $T=2449920 1269520 1 180 $X=2438700 $Y=1269118
X1469 13246 13241 7760 1 3 XNOR2X4 $T=2486880 1229200 1 180 $X=2475660 $Y=1228798
X1470 1745 1 75 1700 3 74 OAI21X4 $T=704880 1309840 0 180 $X=697620 $Y=1304400
X1471 2898 1 2978 2948 3 2893 OAI21X4 $T=893640 1309840 1 180 $X=886380 $Y=1309438
X1472 2841 1 2954 2946 3 3021 OAI21X4 $T=896940 1259440 0 0 $X=896938 $Y=1259038
X1473 2955 1 3023 3015 3 3019 OAI21X4 $T=904200 1360240 1 180 $X=896940 $Y=1359838
X1474 3087 1 3156 3022 3 3158 OAI21X4 $T=924660 1330000 1 180 $X=917400 $Y=1329598
X1475 3357 1 3296 3273 3 3276 OAI21X4 $T=949740 1249360 0 180 $X=942480 $Y=1243920
X1476 3297 1 3356 3374 3 3371 OAI21X4 $T=951720 1289680 0 0 $X=951718 $Y=1289278
X1477 3495 1 3467 3481 3 3420 OAI21X4 $T=980100 1370320 1 180 $X=972840 $Y=1369918
X1478 3735 1 3740 3771 3 156 OAI21X4 $T=1010460 1219120 1 0 $X=1010458 $Y=1213680
X1479 3855 1 3802 3778 3 3708 OAI21X4 $T=1024320 1360240 1 180 $X=1017060 $Y=1359838
X1480 6429 1 6423 6437 3 311 OAI21X4 $T=1430220 1198960 0 0 $X=1430218 $Y=1198558
X1481 6434 1 6339 6379 3 6439 OAI21X4 $T=1437480 1400560 1 180 $X=1430220 $Y=1400158
X1482 6485 1 6506 6630 3 6656 OAI21X4 $T=1461900 1380400 1 0 $X=1461898 $Y=1374960
X1483 6598 1 6658 6660 3 6768 OAI21X4 $T=1464540 1249360 0 0 $X=1464538 $Y=1248958
X1484 6803 1 6672 6827 3 6796 OAI21X4 $T=1487640 1319920 0 0 $X=1487638 $Y=1319518
X1485 6946 1 6952 6921 3 333 OAI21X4 $T=1512060 1158640 1 0 $X=1512058 $Y=1153200
X1486 7058 1 6855 7072 3 7071 OAI21X4 $T=1535820 1209040 1 180 $X=1528560 $Y=1208638
X1487 7092 1 329 7073 3 7089 OAI21X4 $T=1536480 1380400 0 180 $X=1529220 $Y=1374960
X1488 7519 1 7522 7377 3 7501 OAI21X4 $T=1599180 1158640 1 180 $X=1591920 $Y=1158238
X1489 7602 1 7329 7520 3 7708 OAI21X4 $T=1607100 1299760 1 0 $X=1607098 $Y=1294320
X1490 7650 1 7598 7625 3 7686 OAI21X4 $T=1622940 1249360 0 180 $X=1615680 $Y=1243920
X1491 7869 1 7960 7917 3 7959 OAI21X4 $T=1657920 1219120 1 0 $X=1657918 $Y=1213680
X1492 7952 1 7956 7987 3 8091 OAI21X4 $T=1676400 1188880 0 0 $X=1676398 $Y=1188478
X1493 8788 1 8785 8728 3 8764 OAI21X4 $T=1795860 1198960 1 180 $X=1788600 $Y=1198558
X1494 9002 1 8945 8981 3 9003 OAI21X4 $T=1828200 1380400 0 180 $X=1820940 $Y=1374960
X1495 9985 1 9792 10005 3 10010 OAI21X4 $T=1980000 1340080 0 0 $X=1979998 $Y=1339678
X1496 10174 1 10009 10176 3 10077 OAI21X4 $T=2005080 1299760 1 0 $X=2005078 $Y=1294320
X1497 10009 1 10203 10207 3 10231 OAI21X4 $T=2009700 1309840 0 0 $X=2009698 $Y=1309438
X1498 11709 1 11596 11620 3 11707 OAI21X4 $T=2254560 1340080 0 180 $X=2247300 $Y=1334640
X1499 615 1 11875 11853 3 11849 OAI21X4 $T=2288220 1410640 0 0 $X=2288218 $Y=1410238
X1500 11931 1 611 11944 3 11964 OAI21X4 $T=2290860 1370320 0 0 $X=2290858 $Y=1369918
X1501 11960 1 12192 12040 3 12156 OAI21X4 $T=2331780 1309840 0 180 $X=2324520 $Y=1304400
X1502 12040 1 12274 12126 3 12272 OAI21X4 $T=2343660 1289680 1 180 $X=2336400 $Y=1289278
X1503 12463 1 12192 12437 3 12425 OAI21X4 $T=2371380 1299760 0 180 $X=2364120 $Y=1294320
X1504 620 1 12504 12537 3 12540 OAI21X4 $T=2375340 1410640 0 0 $X=2375338 $Y=1410238
X1505 13064 1 12393 13039 3 13038 OAI21X4 $T=2454540 1309840 1 180 $X=2447280 $Y=1309438
X1506 13155 1 13094 13090 3 12992 OAI21X4 $T=2462460 1269520 1 180 $X=2455200 $Y=1269118
X1507 13318 1 13240 13348 3 13347 OAI21X4 $T=2495460 1259440 0 0 $X=2495458 $Y=1259038
X1508 13458 1 13560 13597 3 666 OAI21X4 $T=2518560 1188880 0 0 $X=2518558 $Y=1188478
X1509 14071 1 13941 14059 3 14108 OAI21X4 $T=2589840 1178800 0 0 $X=2589838 $Y=1178398
X1510 4818 1 177 3 CLKBUFX8 $T=1199880 1390480 1 0 $X=1199878 $Y=1385040
X1511 5647 1 295 3 CLKBUFX8 $T=1325280 1279600 1 0 $X=1325278 $Y=1274160
X1512 5648 1 285 3 CLKBUFX8 $T=1327920 1249360 1 0 $X=1327918 $Y=1243920
X1513 8265 1 441 3 CLKBUFX8 $T=1791240 1360240 1 0 $X=1791238 $Y=1354800
X1514 10296 1 10302 3 CLKBUFX8 $T=2026860 1360240 0 0 $X=2026858 $Y=1359838
X1515 12098 1 7393 3 CLKBUFX8 $T=2311320 1340080 0 180 $X=2306700 $Y=1334640
X1516 12901 1 7653 3 CLKBUFX8 $T=2434080 1259440 1 180 $X=2429460 $Y=1259038
X1517 69 1612 3 1 1812 XOR2X2 $T=682440 1330000 1 0 $X=682438 $Y=1324560
X1518 119 3067 3 1 2619 XOR2X2 $T=908820 1138480 1 180 $X=902220 $Y=1138078
X1519 3023 3111 3 1 3423 XOR2X2 $T=910140 1370320 1 0 $X=910138 $Y=1364880
X1520 3467 3466 3 1 2949 XOR2X2 $T=974160 1390480 1 180 $X=967560 $Y=1390078
X1521 3500 142 3 1 139 XOR2X2 $T=979440 1148560 1 180 $X=972840 $Y=1148158
X1522 3703 3695 3 1 153 XOR2X2 $T=1007160 1259440 0 180 $X=1000560 $Y=1254000
X1523 3815 3805 3 1 164 XOR2X2 $T=1026300 1289680 1 180 $X=1019700 $Y=1289278
X1524 4147 4141 3 1 4032 XOR2X2 $T=1073160 1279600 1 180 $X=1066560 $Y=1279198
X1525 101 5465 3 1 266 XOR2X2 $T=1272480 1309840 0 0 $X=1272478 $Y=1309438
X1526 265 5521 3 1 270 XOR2X2 $T=1284360 1350160 0 0 $X=1284358 $Y=1349758
X1527 110 5571 3 1 276 XOR2X2 $T=1290960 1289680 0 0 $X=1290958 $Y=1289278
X1528 104 5576 3 1 280 XOR2X2 $T=1291620 1239280 1 0 $X=1291618 $Y=1233840
X1529 264 5587 3 1 287 XOR2X2 $T=1306800 1350160 1 0 $X=1306798 $Y=1344720
X1530 6457 6482 3 1 6568 XOR2X2 $T=1444740 1289680 1 0 $X=1444738 $Y=1284240
X1531 6658 6661 3 1 6852 XOR2X2 $T=1464540 1269520 1 0 $X=1464538 $Y=1264080
X1532 6724 6506 3 1 7011 XOR2X2 $T=1475100 1380400 1 0 $X=1475098 $Y=1374960
X1533 6762 6769 3 1 6825 XOR2X2 $T=1482360 1229200 0 0 $X=1482358 $Y=1228798
X1534 6877 6947 3 1 7352 XOR2X2 $T=1509420 1168720 0 0 $X=1509418 $Y=1168318
X1535 7179 7172 3 1 7258 XOR2X2 $T=1545720 1249360 1 0 $X=1545718 $Y=1243920
X1536 7421 7443 3 1 7600 XOR2X2 $T=1581360 1188880 1 0 $X=1581358 $Y=1183440
X1537 8759 8752 3 1 439 XOR2X2 $T=1789260 1219120 1 0 $X=1789258 $Y=1213680
X1538 8890 8883 3 1 442 XOR2X2 $T=1808400 1198960 0 180 $X=1801800 $Y=1193520
X1539 8915 8940 3 1 452 XOR2X2 $T=1813020 1198960 1 0 $X=1813018 $Y=1193520
X1540 9952 9947 3 1 9978 XOR2X2 $T=1972080 1330000 0 0 $X=1972078 $Y=1329598
X1541 519 9895 3 1 531 XOR2X2 $T=1972080 1410640 0 0 $X=1972078 $Y=1410238
X1542 10142 10077 3 1 9883 XOR2X2 $T=2001780 1299760 0 180 $X=1995180 $Y=1294320
X1543 518 520 3 1 553 XOR2X2 $T=2035440 1390480 1 0 $X=2035438 $Y=1385040
X1544 12074 12070 3 1 12038 XOR2X2 $T=2310660 1360240 0 180 $X=2304060 $Y=1354800
X1545 12154 12156 3 1 623 XOR2X2 $T=2319900 1309840 0 0 $X=2319898 $Y=1309438
X1546 12245 12244 3 1 12043 XOR2X2 $T=2340360 1410640 1 180 $X=2333760 $Y=1410238
X1547 12293 12287 3 1 12098 XOR2X2 $T=2347620 1340080 0 180 $X=2341020 $Y=1334640
X1548 12280 12192 3 1 627 XOR2X2 $T=2342340 1309840 0 0 $X=2342338 $Y=1309438
X1549 12322 12320 3 1 12132 XOR2X2 $T=2350260 1390480 1 180 $X=2343660 $Y=1390078
X1550 12472 12602 3 1 12650 XOR2X2 $T=2390520 1259440 0 0 $X=2390518 $Y=1259038
X1551 13270 13244 3 1 13129 XOR2X2 $T=2487540 1340080 0 180 $X=2480940 $Y=1334640
X1552 13457 13430 3 1 658 XOR2X2 $T=2507340 1168720 1 180 $X=2500740 $Y=1168318
X1553 13551 13548 3 1 13319 XOR2X2 $T=2519880 1309840 0 180 $X=2513280 $Y=1304400
X1554 13907 13911 3 1 13701 XOR2X2 $T=2564760 1249360 0 180 $X=2558160 $Y=1243920
X1555 14046 13941 3 1 13929 XOR2X2 $T=2582580 1209040 0 180 $X=2575980 $Y=1203600
X1556 67 1 1664 3 INVX2 $T=691020 1259440 0 0 $X=691018 $Y=1259038
X1557 2844 1 2941 3 INVX2 $T=877140 1198960 0 0 $X=877138 $Y=1198558
X1558 2956 1 3065 3 INVX2 $T=894300 1400560 1 0 $X=894298 $Y=1395120
X1559 3019 1 3156 3 INVX2 $T=920040 1350160 1 0 $X=920038 $Y=1344720
X1560 192 1 218 3 INVX2 $T=1152360 1168720 1 180 $X=1150380 $Y=1168318
X1561 4812 1 4451 3 INVX2 $T=1188660 1430800 0 180 $X=1186680 $Y=1425360
X1562 6944 1 6973 3 INVX2 $T=1512060 1390480 0 0 $X=1512058 $Y=1390078
X1563 7543 1 7549 3 INVX2 $T=1597860 1309840 0 0 $X=1597858 $Y=1309438
X1564 7071 1 7632 3 INVX2 $T=1620960 1188880 0 0 $X=1620958 $Y=1188478
X1565 7797 1 7875 3 INVX2 $T=1647360 1219120 0 0 $X=1647358 $Y=1218718
X1566 9665 1 9721 3 INVX2 $T=1935120 1340080 1 0 $X=1935118 $Y=1334640
X1567 9732 1 9689 3 INVX2 $T=1937760 1330000 0 0 $X=1937758 $Y=1329598
X1568 524 1 9703 3 INVX2 $T=1962840 1319920 0 180 $X=1960860 $Y=1314480
X1569 449 1 9853 3 INVX2 $T=1961520 1239280 0 0 $X=1961518 $Y=1238878
X1570 10170 1 10147 3 INVX2 $T=2007720 1269520 1 180 $X=2005740 $Y=1269118
X1571 9930 1 11254 3 INVX2 $T=2187240 1188880 0 0 $X=2187238 $Y=1188478
X1572 13156 1 13096 3 INVX2 $T=2468400 1360240 1 0 $X=2468398 $Y=1354800
X1573 1605 3 1 1655 INVXL $T=693000 1219120 0 0 $X=692998 $Y=1218718
X1574 1917 3 1 1817 INVXL $T=728640 1410640 1 180 $X=727320 $Y=1410238
X1575 1918 3 1 1815 INVXL $T=728640 1420720 1 180 $X=727320 $Y=1420318
X1576 1806 3 1 1942 INVXL $T=731940 1269520 0 0 $X=731938 $Y=1269118
X1577 83 3 1 1842 INVXL $T=737220 1430800 1 0 $X=737218 $Y=1425360
X1578 1980 3 1 1881 INVXL $T=738540 1380400 0 180 $X=737220 $Y=1374960
X1579 2047 3 1 1887 INVXL $T=751740 1380400 1 180 $X=750420 $Y=1379998
X1580 169 3 1 3734 INVXL $T=1036860 1148560 1 180 $X=1035540 $Y=1148158
X1581 221 3 1 4814 INVXL $T=1191300 1380400 0 180 $X=1189980 $Y=1374960
X1582 7406 3 1 7349 INVXL $T=1573440 1249360 1 180 $X=1572120 $Y=1248958
X1583 7466 3 1 7503 INVXL $T=1588620 1400560 1 180 $X=1587300 $Y=1400158
X1584 7839 3 1 7802 INVXL $T=1644720 1269520 1 0 $X=1644718 $Y=1264080
X1585 8887 3 1 8886 INVXL $T=1803120 1188880 0 180 $X=1801800 $Y=1183440
X1586 451 3 1 8859 INVXL $T=1815000 1380400 1 0 $X=1814998 $Y=1374960
X1587 9189 3 1 9209 INVXL $T=1854600 1380400 0 0 $X=1854598 $Y=1379998
X1588 545 3 1 10275 INVXL $T=2036100 1148560 1 180 $X=2034780 $Y=1148158
X1589 10392 3 1 10617 INVXL $T=2079000 1319920 0 0 $X=2078998 $Y=1319518
X1590 11579 3 1 11588 INVXL $T=2238720 1400560 0 0 $X=2238718 $Y=1400158
X1591 12396 3 1 12424 INVXL $T=2361480 1239280 1 0 $X=2361478 $Y=1233840
X1592 645 3 1 13092 INVXL $T=2466420 1420720 1 180 $X=2465100 $Y=1420318
X1593 644 3 1 13183 INVXL $T=2474340 1420720 0 0 $X=2474338 $Y=1420318
X1594 13950 3 1 14050 INVXL $T=2582580 1148560 1 180 $X=2581260 $Y=1148158
X1595 13985 3 1 14076 INVXL $T=2586540 1148560 1 0 $X=2586538 $Y=1143120
X1596 1775 1774 3 1 73 XNOR2X2 $T=707520 1410640 1 180 $X=700260 $Y=1410238
X1597 1751 1773 3 1 84 XNOR2X2 $T=703560 1209040 1 0 $X=703558 $Y=1203600
X1598 1924 1919 3 1 78 XNOR2X2 $T=731280 1390480 0 180 $X=724020 $Y=1385040
X1599 3092 117 3 1 2869 XNOR2X2 $T=911460 1188880 1 180 $X=904200 $Y=1188478
X1600 3110 3113 3 1 2671 XNOR2X2 $T=914100 1168720 1 180 $X=906840 $Y=1168318
X1601 3215 3216 3 1 2917 XNOR2X2 $T=934560 1299760 0 180 $X=927300 $Y=1294320
X1602 3285 3276 3 1 2875 XNOR2X2 $T=948420 1239280 1 180 $X=941160 $Y=1238878
X1603 3351 3296 3 1 2947 XNOR2X2 $T=953700 1269520 0 180 $X=946440 $Y=1264080
X1604 3589 3585 3 1 3550 XNOR2X2 $T=995280 1158640 0 180 $X=988020 $Y=1153200
X1605 3610 3595 3 1 147 XNOR2X2 $T=997920 1188880 0 180 $X=990660 $Y=1183440
X1606 3702 3697 3 1 152 XNOR2X2 $T=1007820 1239280 0 180 $X=1000560 $Y=1233840
X1607 3777 3673 3 1 157 XNOR2X2 $T=1019040 1340080 0 180 $X=1011780 $Y=1334640
X1608 5353 5413 3 1 5488 XNOR2X2 $T=1263900 1168720 1 0 $X=1263898 $Y=1163280
X1609 6399 6406 3 1 6570 XNOR2X2 $T=1428900 1219120 0 0 $X=1428898 $Y=1218718
X1610 6640 6656 3 1 6839 XNOR2X2 $T=1465200 1350160 0 0 $X=1465198 $Y=1349758
X1611 6837 6838 3 1 7010 XNOR2X2 $T=1492920 1219120 1 0 $X=1492918 $Y=1213680
X1612 6802 6868 3 1 6922 XNOR2X2 $T=1497540 1299760 0 0 $X=1497538 $Y=1299358
X1613 6870 6879 3 1 7009 XNOR2X2 $T=1498200 1158640 0 0 $X=1498198 $Y=1158238
X1614 7066 7094 3 1 7264 XNOR2X2 $T=1535160 1138480 0 0 $X=1535158 $Y=1138078
X1615 8073 8091 3 1 8187 XNOR2X2 $T=1680360 1178800 1 0 $X=1680358 $Y=1173360
X1616 429 430 3 1 437 XNOR2X2 $T=1782660 1148560 0 0 $X=1782658 $Y=1148158
X1617 8755 8754 3 1 428 XNOR2X2 $T=1790580 1269520 1 180 $X=1783320 $Y=1269118
X1618 479 9900 3 1 9930 XNOR2X2 $T=1962840 1400560 0 0 $X=1962838 $Y=1400158
X1619 9957 9958 3 1 9855 XNOR2X2 $T=1976040 1309840 0 180 $X=1968780 $Y=1304400
X1620 550 552 3 1 10520 XNOR2X2 $T=2055240 1400560 0 0 $X=2055238 $Y=1400158
X1621 604 9851 3 1 11360 XNOR2X2 $T=2195820 1209040 1 0 $X=2195818 $Y=1203600
X1622 11556 11578 3 1 612 XNOR2X2 $T=2236080 1370320 0 0 $X=2236078 $Y=1369918
X1623 631 632 3 1 12493 XNOR2X2 $T=2366760 1148560 1 0 $X=2366758 $Y=1143120
X1624 12324 12649 3 1 12722 XNOR2X2 $T=2397120 1148560 0 0 $X=2397118 $Y=1148158
X1625 12744 12724 3 1 12502 XNOR2X2 $T=2406360 1360240 0 180 $X=2399100 $Y=1354800
X1626 12743 12802 3 1 12939 XNOR2X2 $T=2432760 1239280 0 0 $X=2432758 $Y=1238878
X1627 13650 13508 3 1 13188 XNOR2X2 $T=2530440 1289680 1 180 $X=2523180 $Y=1289278
X1628 13823 13807 3 1 13561 XNOR2X2 $T=2550240 1269520 0 180 $X=2542980 $Y=1264080
X1629 1610 1607 1 3 42 XOR2X1 $T=685080 1370320 0 180 $X=679800 $Y=1364880
X1630 1633 1631 1 3 63 XOR2X1 $T=691020 1340080 1 180 $X=685740 $Y=1339678
X1631 130 128 1 3 3266 XOR2X1 $T=958980 1209040 1 180 $X=953700 $Y=1208638
X1632 3407 134 1 3 129 XOR2X1 $T=962940 1168720 1 180 $X=957660 $Y=1168318
X1633 3415 136 1 3 131 XOR2X1 $T=964260 1188880 0 180 $X=958980 $Y=1183440
X1634 3464 138 1 3 3349 XOR2X1 $T=972180 1209040 1 180 $X=966900 $Y=1208638
X1635 3867 3864 1 3 168 XOR2X1 $T=1034880 1380400 1 180 $X=1029600 $Y=1379998
X1636 4025 4026 1 3 3796 XOR2X1 $T=1053360 1188880 0 180 $X=1048080 $Y=1183440
X1637 4060 4086 1 3 4025 XOR2X1 $T=1061280 1188880 0 180 $X=1056000 $Y=1183440
X1638 4149 4209 1 3 4147 XOR2X1 $T=1085040 1279600 1 180 $X=1079760 $Y=1279198
X1639 4433 4410 1 3 4117 XOR2X1 $T=1126620 1330000 1 180 $X=1121340 $Y=1329598
X1640 4460 4367 1 3 4433 XOR2X1 $T=1134540 1330000 1 180 $X=1129260 $Y=1329598
X1641 4957 4986 1 3 5061 XOR2X1 $T=1205820 1158640 1 0 $X=1205818 $Y=1153200
X1642 5072 199 1 3 5032 XOR2X1 $T=1221660 1168720 0 180 $X=1216380 $Y=1163280
X1643 5072 4844 1 3 5303 XOR2X1 $T=1222980 1209040 1 0 $X=1222978 $Y=1203600
X1644 5063 5138 1 3 5191 XOR2X1 $T=1228920 1198960 0 0 $X=1228918 $Y=1198558
X1645 250 177 1 3 5262 XOR2X1 $T=1229580 1168720 1 0 $X=1229578 $Y=1163280
X1646 97 5555 1 3 5648 XOR2X1 $T=1296240 1319920 0 0 $X=1296238 $Y=1319518
X1647 274 275 1 3 5647 XOR2X1 $T=1296240 1370320 0 0 $X=1296238 $Y=1369918
X1648 5792 5757 1 3 5810 XOR2X1 $T=1335840 1319920 1 0 $X=1335838 $Y=1314480
X1649 6099 6104 1 3 6342 XOR2X1 $T=1389300 1340080 1 0 $X=1389298 $Y=1334640
X1650 6255 6310 1 3 6671 XOR2X1 $T=1409760 1299760 0 0 $X=1409758 $Y=1299358
X1651 318 316 1 3 6695 XOR2X1 $T=1455960 1138480 0 0 $X=1455958 $Y=1138078
X1652 6659 6704 1 3 6941 XOR2X1 $T=1474440 1400560 1 0 $X=1474438 $Y=1395120
X1653 6975 6972 1 3 7180 XOR2X1 $T=1512060 1330000 0 0 $X=1512058 $Y=1329598
X1654 331 6998 1 3 6696 XOR2X1 $T=1518660 1279600 0 180 $X=1513380 $Y=1274160
X1655 7036 7032 1 3 7005 XOR2X1 $T=1527900 1269520 0 180 $X=1522620 $Y=1264080
X1656 335 7161 1 3 7000 XOR2X1 $T=1545060 1269520 1 180 $X=1539780 $Y=1269118
X1657 7265 7259 1 3 7284 XOR2X1 $T=1555620 1289680 1 0 $X=1555618 $Y=1284240
X1658 7262 7037 1 3 7295 XOR2X1 $T=1555620 1400560 0 0 $X=1555618 $Y=1400158
X1659 7289 7263 1 3 7176 XOR2X1 $T=1560900 1249360 0 180 $X=1555620 $Y=1243920
X1660 7326 7266 1 3 7512 XOR2X1 $T=1563540 1380400 0 0 $X=1563538 $Y=1379998
X1661 340 7376 1 3 341 XOR2X1 $T=1572120 1148560 1 0 $X=1572118 $Y=1143120
X1662 7603 7646 1 3 7792 XOR2X1 $T=1613040 1309840 1 0 $X=1613038 $Y=1304400
X1663 7698 7677 1 3 7921 XOR2X1 $T=1620960 1269520 0 0 $X=1620958 $Y=1269118
X1664 7826 7933 1 3 8098 XOR2X1 $T=1657260 1229200 1 0 $X=1657258 $Y=1223760
X1665 8045 7956 1 3 8117 XOR2X1 $T=1675740 1209040 1 0 $X=1675738 $Y=1203600
X1666 8150 8305 1 3 388 XOR2X1 $T=1710060 1360240 0 0 $X=1710058 $Y=1359838
X1667 8858 8859 1 3 426 XOR2X1 $T=1800480 1380400 0 180 $X=1795200 $Y=1374960
X1668 9075 9074 1 3 459 XOR2X1 $T=1840740 1158640 1 180 $X=1835460 $Y=1158238
X1669 9360 9361 1 3 9245 XOR2X1 $T=1886280 1390480 0 180 $X=1881000 $Y=1385040
X1670 9713 9703 1 3 9664 XOR2X1 $T=1937100 1319920 0 180 $X=1931820 $Y=1314480
X1671 10011 10009 1 3 9923 XOR2X1 $T=1987260 1259440 1 180 $X=1981980 $Y=1259038
X1672 534 10232 1 3 8152 XOR2X1 $T=2016960 1360240 0 180 $X=2011680 $Y=1354800
X1673 548 10387 1 3 10521 XOR2X1 $T=2049960 1420720 1 0 $X=2049958 $Y=1415280
X1674 10767 10768 1 3 575 XOR2X1 $T=2104740 1400560 1 180 $X=2099460 $Y=1400158
X1675 10894 10891 1 3 585 XOR2X1 $T=2128500 1430800 0 180 $X=2123220 $Y=1425360
X1676 11302 11303 1 3 606 XOR2X1 $T=2197140 1370320 0 0 $X=2197138 $Y=1369918
X1677 11791 11811 1 3 12154 XOR2X1 $T=2325840 1299760 0 180 $X=2320560 $Y=1294320
X1678 12568 634 1 3 12870 XOR2X1 $T=2388540 1168720 0 0 $X=2388538 $Y=1168318
X1679 12633 12632 1 3 12434 XOR2X1 $T=2398440 1370320 1 180 $X=2393160 $Y=1369918
X1680 13095 13096 1 3 12957 XOR2X1 $T=2459820 1350160 0 180 $X=2454540 $Y=1344720
X1681 13434 13433 1 3 13420 XOR2X1 $T=2507340 1400560 0 180 $X=2502060 $Y=1395120
X1682 663 13525 1 3 13519 XOR2X1 $T=2520540 1400560 0 180 $X=2515260 $Y=1395120
X1683 13696 13219 1 3 13680 XOR2X1 $T=2537700 1380400 0 180 $X=2532420 $Y=1374960
X1684 13805 13815 1 3 13875 XOR2X1 $T=2546940 1390480 0 0 $X=2546938 $Y=1390078
X1685 14078 14072 1 3 13881 XOR2X1 $T=2586540 1229200 1 180 $X=2581260 $Y=1228798
X1686 14336 14335 1 3 14313 XOR2X1 $T=2622840 1360240 1 180 $X=2617560 $Y=1359838
X1687 1549 3 1605 1606 1 NOR2BX1 $T=689700 1249360 0 180 $X=687060 $Y=1243920
X1688 2167 3 2113 1610 1 NOR2BX1 $T=756360 1370320 1 180 $X=753720 $Y=1369918
X1689 3273 3 3357 3351 1 NOR2BX1 $T=956340 1249360 1 180 $X=953700 $Y=1248958
X1690 3478 3 3434 3405 1 NOR2BX1 $T=977460 1309840 1 180 $X=974820 $Y=1309438
X1691 156 3 3671 3675 1 NOR2BX1 $T=1010460 1178800 0 0 $X=1010458 $Y=1178398
X1692 3711 3 3694 3610 1 NOR2BX1 $T=1020360 1168720 1 180 $X=1017720 $Y=1168318
X1693 4669 3 4666 4665 1 NOR2BX1 $T=1162920 1198960 0 180 $X=1160280 $Y=1193520
X1694 5019 3 5022 5185 1 NOR2BX1 $T=1228260 1229200 1 0 $X=1228258 $Y=1223760
X1695 8862 3 8882 8915 1 NOR2BX1 $T=1813020 1168720 1 180 $X=1810380 $Y=1168318
X1696 9960 3 9959 9952 1 NOR2BX1 $T=1976700 1360240 0 180 $X=1974060 $Y=1354800
X1697 11526 3 11546 11556 1 NOR2BX1 $T=2231460 1360240 1 0 $X=2231458 $Y=1354800
X1698 12328 3 12397 12323 1 NOR2BX1 $T=2360820 1420720 0 180 $X=2358180 $Y=1415280
X1699 661 3 660 13434 1 NOR2BX1 $T=2507340 1410640 0 180 $X=2504700 $Y=1405200
X1700 13317 3 13287 13418 1 NOR2BX1 $T=2512620 1198960 1 180 $X=2509980 $Y=1198558
X1701 654 3 660 13552 1 NOR2BX1 $T=2515260 1420720 0 0 $X=2515258 $Y=1420318
X1702 14082 3 14064 14138 1 NOR2BX1 $T=2599080 1158640 1 180 $X=2596440 $Y=1158238
X1703 102 2339 2303 2245 3 1 2182 ADDFX2 $T=790680 1420720 1 180 $X=776820 $Y=1420318
X1704 2515 2383 2354 2242 3 1 2232 ADDFX2 $T=799920 1330000 1 180 $X=786060 $Y=1329598
X1705 91 95 2399 2380 3 1 2341 ADDFX2 $T=806520 1209040 1 180 $X=792660 $Y=1208638
X1706 2463 2469 2464 2307 3 1 2208 ADDFX2 $T=811800 1400560 1 180 $X=797940 $Y=1400158
X1707 2545 2490 96 2463 3 1 2303 ADDFX2 $T=811800 1420720 0 180 $X=797940 $Y=1415280
X1708 2524 2512 2485 2330 3 1 2370 ADDFX2 $T=814440 1239280 1 180 $X=800580 $Y=1238878
X1709 2468 2516 2467 2336 3 1 2282 ADDFX2 $T=815100 1380400 0 180 $X=801240 $Y=1374960
X1710 2544 2517 2489 2467 3 1 2464 ADDFX2 $T=815760 1390480 1 180 $X=801900 $Y=1390078
X1711 2542 2521 2491 2371 3 1 2309 ADDFX2 $T=817080 1299760 1 180 $X=803220 $Y=1299358
X1712 2567 98 2487 2486 3 1 2468 ADDFX2 $T=817740 1380400 1 180 $X=803880 $Y=1379998
X1713 2486 2488 2493 2236 3 1 2342 ADDFX2 $T=818400 1340080 1 180 $X=804540 $Y=1339678
X1714 99 100 2512 2383 3 1 2488 ADDFX2 $T=819720 1319920 0 180 $X=805860 $Y=1314480
X1715 105 87 2522 2515 3 1 2493 ADDFX2 $T=822360 1350160 1 180 $X=808500 $Y=1349758
X1716 97 104 2523 2491 3 1 2354 ADDFX2 $T=823020 1330000 0 180 $X=809160 $Y=1324560
X1717 2589 103 2514 2374 3 1 2518 ADDFX2 $T=825000 1249360 1 180 $X=811140 $Y=1248958
X1718 100 2512 107 2573 3 1 2542 ADDFX2 $T=813780 1309840 0 0 $X=813778 $Y=1309438
X1719 95 99 108 2589 3 1 2549 ADDFX2 $T=814440 1269520 1 0 $X=814438 $Y=1264080
X1720 2573 109 2549 2543 3 1 2404 ADDFX2 $T=828960 1279600 1 180 $X=815100 $Y=1279198
X1721 4279 4145 4117 4022 3 1 3877 ADDFX2 $T=1075800 1330000 1 180 $X=1061940 $Y=1329598
X1722 4280 4191 4178 4021 3 1 4093 ADDFX2 $T=1085040 1360240 1 180 $X=1071180 $Y=1359838
X1723 4343 4204 4182 3841 3 1 3905 ADDFX2 $T=1086360 1209040 1 180 $X=1072500 $Y=1208638
X1724 4241 177 4183 4089 3 1 4146 ADDFX2 $T=1086360 1380400 0 180 $X=1072500 $Y=1374960
X1725 4247 179 4188 176 3 1 4060 ADDFX2 $T=1089000 1168720 1 180 $X=1075140 $Y=1168318
X1726 4263 4240 4206 4086 3 1 4182 ADDFX2 $T=1091640 1198960 1 180 $X=1077780 $Y=1198558
X1727 4339 4246 181 178 3 1 3904 ADDFX2 $T=1094940 1148560 1 180 $X=1081080 $Y=1148158
X1728 180 177 4269 4273 3 1 4345 ADDFX2 $T=1084380 1249360 0 0 $X=1084378 $Y=1248958
X1729 4340 180 4273 4206 3 1 4143 ADDFX2 $T=1103520 1229200 1 180 $X=1089660 $Y=1228798
X1730 187 185 4269 4149 3 1 4264 ADDFX2 $T=1104840 1289680 1 180 $X=1090980 $Y=1289278
X1731 184 179 182 4188 3 1 4240 ADDFX2 $T=1106160 1178800 0 180 $X=1092300 $Y=1173360
X1732 187 4307 4303 4266 3 1 4186 ADDFX2 $T=1107480 1390480 1 180 $X=1093620 $Y=1390078
X1733 196 192 4306 4279 3 1 4125 ADDFX2 $T=1108140 1340080 1 180 $X=1094280 $Y=1339678
X1734 191 193 4307 4280 3 1 4183 ADDFX2 $T=1108140 1370320 1 180 $X=1094280 $Y=1369918
X1735 198 189 186 4301 3 1 4145 ADDFX2 $T=1109460 1330000 0 180 $X=1095600 $Y=1324560
X1736 183 177 186 4205 3 1 4178 ADDFX2 $T=1110120 1360240 0 180 $X=1096260 $Y=1354800
X1737 4409 4363 4342 4339 3 1 4026 ADDFX2 $T=1112760 1168720 1 180 $X=1098900 $Y=1168318
X1738 189 194 4367 4366 3 1 4392 ADDFX2 $T=1101540 1279600 0 0 $X=1101538 $Y=1279198
X1739 4437 197 4346 4342 3 1 4204 ADDFX2 $T=1115400 1198960 1 180 $X=1101540 $Y=1198558
X1740 4430 4369 4347 4343 3 1 4062 ADDFX2 $T=1115400 1219120 1 180 $X=1101540 $Y=1218718
X1741 4345 4366 4361 4095 3 1 4457 ADDFX2 $T=1104840 1249360 0 0 $X=1104838 $Y=1248958
X1742 4426 200 4368 195 3 1 4246 ADDFX2 $T=1120020 1148560 1 180 $X=1106160 $Y=1148158
X1743 199 194 4383 4347 3 1 4361 ADDFX2 $T=1120680 1239280 1 180 $X=1106820 $Y=1238878
X1744 177 183 199 4247 3 1 4263 ADDFX2 $T=1122000 1209040 0 180 $X=1108140 $Y=1203600
X1745 192 193 204 4426 3 1 4409 ADDFX2 $T=1135860 1168720 0 180 $X=1122000 $Y=1163280
X1746 192 197 204 4346 3 1 4369 ADDFX2 $T=1139160 1198960 0 180 $X=1125300 $Y=1193520
X1747 205 191 4459 4437 3 1 4430 ADDFX2 $T=1139160 1219120 0 180 $X=1125300 $Y=1213680
X1748 185 200 208 4368 3 1 4363 ADDFX2 $T=1143780 1148560 1 180 $X=1129920 $Y=1148158
X1749 205 209 4459 4511 3 1 4484 ADDFX2 $T=1130580 1229200 1 0 $X=1130578 $Y=1223760
X1750 196 209 210 4479 3 1 4214 ADDFX2 $T=1144440 1309840 0 180 $X=1130580 $Y=1304400
X1751 193 184 210 4410 3 1 4157 ADDFX2 $T=1144440 1340080 0 180 $X=1130580 $Y=1334640
X1752 5835 288 295 5996 3 1 6027 ADDFX2 $T=1356300 1239280 1 0 $X=1356298 $Y=1233840
X1753 294 290 6027 6044 3 1 6135 ADDFX2 $T=1362240 1259440 0 0 $X=1362238 $Y=1259038
X1754 5973 290 6036 6046 3 1 6000 ADDFX2 $T=1362900 1309840 1 0 $X=1362898 $Y=1304400
X1755 5996 287 6132 6149 3 1 6253 ADDFX2 $T=1379400 1229200 0 0 $X=1379398 $Y=1228798
X1756 295 5973 299 6103 3 1 6132 ADDFX2 $T=1380720 1239280 1 0 $X=1380718 $Y=1233840
X1757 295 296 299 301 3 1 6156 ADDFX2 $T=1382700 1148560 0 0 $X=1382698 $Y=1148158
X1758 270 5945 6156 6164 3 1 6157 ADDFX2 $T=1384020 1168720 1 0 $X=1384018 $Y=1163280
X1759 294 287 5946 6127 3 1 6158 ADDFX2 $T=1384020 1209040 1 0 $X=1384018 $Y=1203600
X1760 6103 270 6158 6165 3 1 6251 ADDFX2 $T=1384020 1219120 1 0 $X=1384018 $Y=1213680
X1761 299 5973 294 6191 3 1 6257 ADDFX2 $T=1387320 1279600 0 0 $X=1387318 $Y=1279198
X1762 10628 10478 10431 10266 3 1 10297 ADDFX2 $T=2058540 1209040 1 180 $X=2044680 $Y=1208638
X1763 10475 10498 10479 10431 3 1 10299 ADDFX2 $T=2062500 1229200 1 180 $X=2048640 $Y=1228798
X1764 10529 554 549 10478 3 1 10475 ADDFX2 $T=2064480 1239280 0 180 $X=2050620 $Y=1233840
X1765 10601 549 10526 10479 3 1 10480 ADDFX2 $T=2073720 1249360 1 180 $X=2059860 $Y=1248958
X1766 555 558 10553 10526 3 1 10531 ADDFX2 $T=2061180 1279600 0 0 $X=2061178 $Y=1279198
X1767 10529 558 567 10619 3 1 10628 ADDFX2 $T=2071740 1198960 0 0 $X=2071738 $Y=1198558
X1768 570 568 10575 10322 3 1 10432 ADDFX2 $T=2085600 1148560 1 180 $X=2071740 $Y=1148158
X1769 560 10579 10576 561 3 1 10496 ADDFX2 $T=2085600 1168720 1 180 $X=2071740 $Y=1168318
X1770 10619 560 10569 10575 3 1 10238 ADDFX2 $T=2085600 1178800 0 180 $X=2071740 $Y=1173360
X1771 567 10601 563 10576 3 1 10569 ADDFX2 $T=2085600 1188880 0 180 $X=2071740 $Y=1183440
X1772 549 10572 10498 10585 3 1 10579 ADDFX2 $T=2087580 1229200 1 180 $X=2073720 $Y=1228798
X1773 10558 10529 10585 565 3 1 564 ADDFX2 $T=2089560 1209040 0 180 $X=2075700 $Y=1203600
X1774 573 567 10766 576 3 1 574 ADDFX2 $T=2113980 1148560 0 180 $X=2100120 $Y=1143120
X1775 555 10815 10553 577 3 1 10766 ADDFX2 $T=2114640 1229200 1 180 $X=2100780 $Y=1228798
X1776 10769 9930 10819 580 3 1 583 ADDFX2 $T=2104080 1168720 0 0 $X=2104078 $Y=1168318
X1777 573 549 10814 10783 3 1 578 ADDFX2 $T=2118600 1158640 1 180 $X=2104740 $Y=1158238
X1778 570 10783 559 10819 3 1 582 ADDFX2 $T=2105400 1158640 1 0 $X=2105398 $Y=1153200
X1779 10529 567 10862 10866 3 1 10823 ADDFX2 $T=2112000 1340080 0 0 $X=2111998 $Y=1339678
X1780 10886 10897 553 589 3 1 590 ADDFX2 $T=2125860 1198960 1 0 $X=2125858 $Y=1193520
X1781 10529 558 549 10940 3 1 10886 ADDFX2 $T=2125860 1198960 0 0 $X=2125858 $Y=1198558
X1782 10956 554 555 10897 3 1 10814 ADDFX2 $T=2140380 1229200 1 180 $X=2126520 $Y=1228798
X1783 560 570 10925 587 3 1 10889 ADDFX2 $T=2144340 1370320 0 180 $X=2130480 $Y=1364880
X1784 10984 10940 559 588 3 1 10769 ADDFX2 $T=2145000 1168720 1 180 $X=2131140 $Y=1168318
X1785 567 560 10941 10893 3 1 10865 ADDFX2 $T=2146980 1340080 1 180 $X=2133120 $Y=1339678
X1786 10925 554 559 11009 3 1 11235 ADDFX2 $T=2135760 1299760 0 0 $X=2135758 $Y=1299358
X1787 10529 555 567 591 3 1 10984 ADDFX2 $T=2156220 1188880 0 180 $X=2142360 $Y=1183440
X1788 567 549 573 594 3 1 595 ADDFX2 $T=2146980 1148560 0 0 $X=2146978 $Y=1148158
X1789 560 10529 553 596 3 1 597 ADDFX2 $T=2150280 1138480 0 0 $X=2150278 $Y=1138078
X1790 11030 10520 11121 11125 3 1 11071 ADDFX2 $T=2153580 1390480 1 0 $X=2153578 $Y=1385040
X1791 11091 11009 551 11148 3 1 11362 ADDFX2 $T=2157540 1289680 1 0 $X=2157538 $Y=1284240
X1792 10302 559 10941 11175 3 1 11176 ADDFX2 $T=2162820 1319920 0 0 $X=2162818 $Y=1319518
X1793 573 553 10862 11126 3 1 11123 ADDFX2 $T=2177340 1340080 0 180 $X=2163480 $Y=1334640
X1794 11126 11150 11176 11182 3 1 11412 ADDFX2 $T=2165460 1330000 0 0 $X=2165458 $Y=1329598
X1795 11147 11250 11123 11285 3 1 11259 ADDFX2 $T=2183940 1350160 0 0 $X=2183938 $Y=1349758
X1796 11235 11175 11275 11356 3 1 11357 ADDFX2 $T=2187900 1299760 0 0 $X=2187898 $Y=1299358
X1797 11390 543 11287 11283 3 1 11275 ADDFX2 $T=2205720 1269520 1 180 $X=2191860 $Y=1269118
X1798 525 567 11390 11447 3 1 11708 ADDFX2 $T=2205060 1249360 0 0 $X=2205058 $Y=1248958
X1799 11538 531 10946 11604 3 1 11606 ADDFX2 $T=2230800 1269520 0 0 $X=2230798 $Y=1269118
X1800 11619 11254 11178 11732 3 1 11733 ADDFX2 $T=2244000 1239280 1 0 $X=2243998 $Y=1233840
X1801 553 609 11598 11752 3 1 11759 ADDFX2 $T=2248620 1158640 1 0 $X=2248618 $Y=1153200
X1802 559 605 11761 11786 3 1 11804 ADDFX2 $T=2255880 1138480 0 0 $X=2255878 $Y=1138078
X1803 11736 525 11785 11787 3 1 11792 ADDFX2 $T=2257200 1259440 0 0 $X=2257198 $Y=1259038
X1804 531 549 11250 11785 3 1 11755 ADDFX2 $T=2257200 1289680 1 0 $X=2257198 $Y=1284240
X1805 11604 11755 11733 11791 3 1 11927 ADDFX2 $T=2257200 1299760 1 0 $X=2257198 $Y=1294320
X1806 10172 614 11619 11818 3 1 11757 ADDFX2 $T=2261820 1188880 0 0 $X=2261818 $Y=1188478
X1807 11757 11614 11639 11821 3 1 11826 ADDFX2 $T=2262480 1198960 1 0 $X=2262478 $Y=1193520
X1808 11814 609 11447 11869 3 1 11934 ADDFX2 $T=2273040 1209040 0 0 $X=2273038 $Y=1208638
X1809 11869 11882 11698 11926 3 1 11962 ADDFX2 $T=2280960 1209040 1 0 $X=2280958 $Y=1203600
X1810 522 11883 11912 11882 3 1 11911 ADDFX2 $T=2280960 1229200 0 0 $X=2280958 $Y=1228798
X1811 573 522 11736 11943 3 1 11969 ADDFX2 $T=2284260 1178800 0 0 $X=2284258 $Y=1178398
X1812 11810 11911 11934 11963 3 1 12165 ADDFX2 $T=2285580 1229200 1 0 $X=2285578 $Y=1223760
X1813 543 608 11786 11965 3 1 12072 ADDFX2 $T=2286240 1138480 0 0 $X=2286238 $Y=1138078
X1814 11969 12042 11818 12131 3 1 12102 ADDFX2 $T=2307360 1188880 0 0 $X=2307358 $Y=1188478
X1815 11943 622 11759 12212 3 1 12220 ADDFX2 $T=2319900 1168720 1 0 $X=2319898 $Y=1163280
X1816 1777 1776 1 3 70 XNOR2X1 $T=708180 1330000 1 180 $X=702900 $Y=1329598
X1817 1993 1986 1 3 80 XNOR2X1 $T=742500 1299760 1 180 $X=737220 $Y=1299358
X1818 87 2107 1 3 1923 XNOR2X1 $T=755040 1178800 0 180 $X=749760 $Y=1173360
X1819 2114 2115 1 3 1541 XNOR2X1 $T=755040 1219120 0 180 $X=749760 $Y=1213680
X1820 2136 2137 1 3 1897 XNOR2X1 $T=757020 1279600 0 180 $X=751740 $Y=1274160
X1821 2158 2157 1 3 1865 XNOR2X1 $T=760980 1289680 1 180 $X=755700 $Y=1289278
X1822 2179 2180 1 3 1601 XNOR2X1 $T=766260 1239280 0 180 $X=760980 $Y=1233840
X1823 2341 2330 1 3 2114 XNOR2X1 $T=802560 1219120 0 180 $X=797280 $Y=1213680
X1824 99 87 1 3 2403 XNOR2X1 $T=815100 1178800 1 180 $X=809820 $Y=1178398
X1825 106 99 1 3 2545 XNOR2X1 $T=823020 1430800 0 180 $X=817740 $Y=1425360
X1826 99 108 1 3 2524 XNOR2X1 $T=825660 1239280 1 180 $X=820380 $Y=1238878
X1827 127 3372 1 3 3114 XNOR2X1 $T=956340 1410640 1 180 $X=951060 $Y=1410238
X1828 3406 3420 1 3 2951 XNOR2X1 $T=964920 1370320 1 180 $X=959640 $Y=1369918
X1829 3741 3732 1 3 155 XNOR2X1 $T=1013760 1289680 0 180 $X=1008480 $Y=1284240
X1830 3834 3816 1 3 163 XNOR2X1 $T=1026960 1380400 1 180 $X=1021680 $Y=1379998
X1831 4053 4051 1 3 170 XNOR2X1 $T=1058640 1410640 0 180 $X=1053360 $Y=1405200
X1832 198 192 1 3 4191 XNOR2X1 $T=1122660 1350160 0 180 $X=1117380 $Y=1344720
X1833 185 184 1 3 4460 XNOR2X1 $T=1137180 1330000 0 0 $X=1137178 $Y=1329598
X1834 198 210 1 3 4807 XNOR2X1 $T=1181400 1249360 0 0 $X=1181398 $Y=1248958
X1835 228 232 1 3 5108 XNOR2X1 $T=1209120 1249360 0 0 $X=1209118 $Y=1248958
X1836 230 191 1 3 5072 XNOR2X1 $T=1215060 1289680 1 0 $X=1215058 $Y=1284240
X1837 5032 5061 1 3 5236 XNOR2X1 $T=1218360 1158640 1 0 $X=1218358 $Y=1153200
X1838 228 188 1 3 5138 XNOR2X1 $T=1218360 1219120 1 0 $X=1218358 $Y=1213680
X1839 5109 249 1 3 5241 XNOR2X1 $T=1228260 1299760 1 0 $X=1228258 $Y=1294320
X1840 4954 187 1 3 250 XNOR2X1 $T=1236180 1178800 0 180 $X=1230900 $Y=1173360
X1841 5264 253 1 3 5413 XNOR2X1 $T=1254660 1168720 0 0 $X=1254658 $Y=1168318
X1842 235 5585 1 3 278 XNOR2X1 $T=1296240 1269520 0 0 $X=1296238 $Y=1269118
X1843 5668 5488 1 3 6004 XNOR2X1 $T=1308120 1158640 0 0 $X=1308118 $Y=1158238
X1844 5553 5487 1 3 5668 XNOR2X1 $T=1313400 1168720 1 180 $X=1308120 $Y=1168318
X1845 5652 5716 1 3 5742 XNOR2X1 $T=1321320 1158640 1 0 $X=1321318 $Y=1153200
X1846 188 247 1 3 5792 XNOR2X1 $T=1327920 1319920 1 0 $X=1327918 $Y=1314480
X1847 186 6105 1 3 300 XNOR2X1 $T=1382700 1360240 1 0 $X=1382698 $Y=1354800
X1848 6260 6283 1 3 6666 XNOR2X1 $T=1407780 1330000 0 0 $X=1407778 $Y=1329598
X1849 6149 6251 1 3 6399 XNOR2X1 $T=1414380 1219120 0 0 $X=1414378 $Y=1218718
X1850 6426 6309 1 3 6595 XNOR2X1 $T=1431540 1249360 0 0 $X=1431538 $Y=1248958
X1851 6569 6505 1 3 6627 XNOR2X1 $T=1451340 1198960 0 0 $X=1451338 $Y=1198558
X1852 6478 6675 1 3 6725 XNOR2X1 $T=1470480 1410640 1 0 $X=1470478 $Y=1405200
X1853 6880 6878 1 3 324 XNOR2X1 $T=1501500 1410640 0 180 $X=1496220 $Y=1405200
X1854 7160 7353 1 3 7472 XNOR2X1 $T=1568820 1360240 0 0 $X=1568818 $Y=1359838
X1855 7395 7390 1 3 7531 XNOR2X1 $T=1576080 1350160 1 0 $X=1576078 $Y=1344720
X1856 342 7388 1 3 7391 XNOR2X1 $T=1581360 1269520 1 180 $X=1576080 $Y=1269118
X1857 344 7348 1 3 346 XNOR2X1 $T=1589280 1229200 0 0 $X=1589278 $Y=1228798
X1858 7647 7622 1 3 7753 XNOR2X1 $T=1613040 1309840 0 0 $X=1613038 $Y=1309438
X1859 7718 7719 1 3 7833 XNOR2X1 $T=1626240 1259440 1 0 $X=1626238 $Y=1254000
X1860 7918 7876 1 3 7962 XNOR2X1 $T=1651980 1239280 1 0 $X=1651978 $Y=1233840
X1861 7989 368 1 3 8007 XNOR2X1 $T=1671780 1380400 0 180 $X=1666500 $Y=1374960
X1862 369 371 1 3 8151 XNOR2X1 $T=1673760 1148560 1 0 $X=1673758 $Y=1143120
X1863 8264 8267 1 3 386 XNOR2X1 $T=1704780 1330000 0 0 $X=1704778 $Y=1329598
X1864 8363 8495 1 3 409 XNOR2X1 $T=1746360 1299760 0 180 $X=1741080 $Y=1294320
X1865 8707 8704 1 3 8684 XNOR2X1 $T=1780680 1229200 1 180 $X=1775400 $Y=1228798
X1866 8889 8865 1 3 8918 XNOR2X1 $T=1806420 1360240 1 0 $X=1806418 $Y=1354800
X1867 8951 8948 1 3 8922 XNOR2X1 $T=1819620 1390480 0 180 $X=1814340 $Y=1385040
X1868 9077 9073 1 3 460 XNOR2X1 $T=1841400 1148560 1 180 $X=1836120 $Y=1148158
X1869 9325 9323 1 3 9240 XNOR2X1 $T=1879680 1410640 0 180 $X=1874400 $Y=1405200
X1870 9628 9627 1 3 9592 XNOR2X1 $T=1923240 1330000 1 180 $X=1917960 $Y=1329598
X1871 10274 10275 1 3 8941 XNOR2X1 $T=2026200 1158640 0 180 $X=2020920 $Y=1153200
X1872 535 10268 1 3 10296 XNOR2X1 $T=2023560 1420720 0 0 $X=2023558 $Y=1420318
X1873 10172 570 1 3 586 XNOR2X1 $T=2136420 1390480 0 180 $X=2131140 $Y=1385040
X1874 11182 11357 1 3 11302 XNOR2X1 $T=2203080 1340080 0 180 $X=2197800 $Y=1334640
X1875 11455 11451 1 3 607 XNOR2X1 $T=2219580 1410640 1 180 $X=2214300 $Y=1410238
X1876 12500 12559 1 3 12628 XNOR2X1 $T=2391180 1269520 1 0 $X=2391178 $Y=1264080
X1877 636 635 1 3 12713 XNOR2X1 $T=2405700 1420720 1 180 $X=2400420 $Y=1420318
X1878 12571 12817 1 3 12844 XNOR2X1 $T=2418900 1239280 0 0 $X=2418898 $Y=1238878
X1879 640 639 1 3 12874 XNOR2X1 $T=2434080 1430800 0 180 $X=2428800 $Y=1425360
X1880 12564 12905 1 3 13093 XNOR2X1 $T=2434080 1219120 0 0 $X=2434078 $Y=1218718
X1881 12935 12956 1 3 13122 XNOR2X1 $T=2439360 1158640 0 0 $X=2439358 $Y=1158238
X1882 12993 12978 1 3 12906 XNOR2X1 $T=2448600 1390480 1 180 $X=2443320 $Y=1390078
X1883 13098 13094 1 3 12901 XNOR2X1 $T=2460480 1259440 1 180 $X=2455200 $Y=1259038
X1884 13181 13180 1 3 13123 XNOR2X1 $T=2473680 1380400 1 180 $X=2468400 $Y=1379998
X1885 13278 13286 1 3 13305 XNOR2X1 $T=2488860 1158640 0 0 $X=2488858 $Y=1158238
X1886 13765 13763 1 3 662 XNOR2X1 $T=2544300 1148560 0 180 $X=2539020 $Y=1143120
X1887 675 13869 1 3 13787 XNOR2X1 $T=2552880 1360240 1 180 $X=2547600 $Y=1359838
X1888 13946 13951 1 3 13966 XNOR2X1 $T=2564760 1400560 0 0 $X=2564758 $Y=1400158
X1889 13986 13981 1 3 13967 XNOR2X1 $T=2572680 1360240 0 180 $X=2567400 $Y=1354800
X1890 687 14017 1 3 14079 XNOR2X1 $T=2577960 1400560 1 0 $X=2577958 $Y=1395120
X1891 688 675 1 3 14110 XNOR2X1 $T=2588520 1380400 0 0 $X=2588518 $Y=1379998
X1892 5347 5260 1 198 3 256 5177 5243 OAI221XL $T=1244100 1390480 1 180 $X=1239480 $Y=1390078
X1893 12369 12292 1 12527 3 12534 12456 12723 OAI221XL $T=2377320 1198960 0 0 $X=2377318 $Y=1198558
X1894 14041 13219 1 13877 3 14009 682 14017 OAI221XL $T=2577960 1410640 0 180 $X=2573340 $Y=1405200
X1895 14280 13219 1 14277 3 14257 14226 14256 OAI221XL $T=2612940 1370320 0 180 $X=2608320 $Y=1364880
X1896 188 4303 183 3 1 4241 ADDHXL $T=1103520 1390480 0 180 $X=1096260 $Y=1385040
X1897 187 4383 188 3 1 4340 ADDHXL $T=1119360 1229200 1 180 $X=1112100 $Y=1228798
X1898 304 6493 303 3 1 6667 ADDHXL $T=1454640 1420720 0 0 $X=1454638 $Y=1420318
X1899 6667 6676 314 3 1 6797 ADDHXL $T=1479060 1420720 0 0 $X=1479058 $Y=1420318
X1900 6797 6974 325 3 1 7450 ADDHXL $T=1508760 1410640 0 0 $X=1508758 $Y=1410238
X1901 7450 7454 7465 3 1 7524 ADDHXL $T=1582680 1410640 1 0 $X=1582678 $Y=1405200
X1902 7517 7550 7526 3 1 7678 ADDHXL $T=1595220 1340080 1 0 $X=1595218 $Y=1334640
X1903 7524 7552 7521 3 1 7551 ADDHXL $T=1595220 1380400 0 0 $X=1595218 $Y=1379998
X1904 7551 7532 7523 3 1 7517 ADDHXL $T=1602480 1370320 0 180 $X=1595220 $Y=1364880
X1905 7796 7829 7838 3 1 7850 ADDHXL $T=1639440 1309840 1 0 $X=1639438 $Y=1304400
X1906 7678 7841 7821 3 1 7796 ADDHXL $T=1650000 1319920 1 180 $X=1642740 $Y=1319518
X1907 7850 7925 7920 3 1 8014 ADDHXL $T=1650000 1279600 1 0 $X=1649998 $Y=1274160
X1908 8014 8036 7924 3 1 8046 ADDHXL $T=1668480 1269520 1 0 $X=1668478 $Y=1264080
X1909 8046 8145 8242 3 1 8297 ADDHXL $T=1694220 1249360 0 0 $X=1694218 $Y=1248958
X1910 8276 8296 8303 3 1 8333 ADDHXL $T=1706100 1168720 1 0 $X=1706098 $Y=1163280
X1911 8297 8304 8311 3 1 8332 ADDHXL $T=1707420 1249360 1 0 $X=1707418 $Y=1243920
X1912 8313 8263 8335 3 1 8339 ADDHXL $T=1712700 1188880 1 0 $X=1712698 $Y=1183440
X1913 8332 8327 8277 3 1 8313 ADDHXL $T=1720620 1229200 0 180 $X=1713360 $Y=1223760
X1914 8333 8274 392 3 1 8397 ADDHXL $T=1715340 1138480 0 0 $X=1715338 $Y=1138078
X1915 8339 8368 8373 3 1 8276 ADDHXL $T=1717320 1168720 0 0 $X=1717318 $Y=1168318
X1916 9098 9070 422 3 1 468 ADDHXL $T=1840740 1400560 1 0 $X=1840738 $Y=1395120
X1917 465 9066 423 3 1 9098 ADDHXL $T=1848660 1420720 0 180 $X=1841400 $Y=1415280
X1918 9590 9572 9504 3 1 9660 ADDHXL $T=1912680 1209040 1 0 $X=1912678 $Y=1203600
X1919 496 9595 9443 3 1 9590 ADDHXL $T=1923900 1158640 1 180 $X=1916640 $Y=1158238
X1920 9620 9596 9328 3 1 9558 ADDHXL $T=1923900 1279600 1 180 $X=1916640 $Y=1279198
X1921 9660 9683 9506 3 1 9724 ADDHXL $T=1927200 1209040 1 0 $X=1927198 $Y=1203600
X1922 9688 9667 9347 3 1 9620 ADDHXL $T=1934460 1259440 0 180 $X=1927200 $Y=1254000
X1923 9725 9710 9386 3 1 9688 ADDHXL $T=1939740 1239280 0 180 $X=1932480 $Y=1233840
X1924 9724 9735 9508 3 1 9725 ADDHXL $T=1935120 1229200 0 0 $X=1935118 $Y=1228798
X1925 555 10601 556 3 1 10498 ADDHXL $T=2082300 1239280 0 180 $X=2075040 $Y=1233840
X1926 554 10572 556 3 1 10676 ADDHXL $T=2090220 1289680 0 0 $X=2090218 $Y=1289278
X1927 558 10815 556 3 1 10956 ADDHXL $T=2111340 1239280 1 0 $X=2111338 $Y=1233840
X1928 553 11150 556 3 1 11287 ADDHXL $T=2168100 1299760 1 0 $X=2168098 $Y=1294320
X1929 3 1748 62 1779 1 NOR2XL $T=705540 1239280 0 0 $X=705538 $Y=1238878
X1930 3 377 370 382 1 NOR2XL $T=1691580 1420720 1 0 $X=1691578 $Y=1415280
X1931 3 556 10497 10394 1 NOR2XL $T=2058540 1360240 0 180 $X=2056560 $Y=1354800
X1932 3 14228 14257 14143 1 NOR2XL $T=2607000 1370320 0 0 $X=2606998 $Y=1369918
X1933 2299 2269 91 1 3 90 XOR3X2 $T=783420 1158640 0 180 $X=771540 $Y=1153200
X1934 2350 2380 2403 1 3 92 XOR3X2 $T=790020 1178800 0 0 $X=790018 $Y=1178398
X1935 134 162 159 1 3 3505 XOR3X2 $T=1023660 1430800 0 180 $X=1011780 $Y=1425360
X1936 4778 208 218 1 3 4986 XOR3X2 $T=1182060 1148560 1 0 $X=1182058 $Y=1143120
X1937 4947 4952 4953 1 3 241 XOR3X2 $T=1201200 1198960 1 0 $X=1201198 $Y=1193520
X1938 5226 204 5303 1 3 5520 XOR3X2 $T=1239480 1188880 0 0 $X=1239478 $Y=1188478
X1939 5435 5354 4811 1 3 5498 XOR3X2 $T=1269180 1229200 0 0 $X=1269178 $Y=1228798
X1940 290 288 5835 1 3 5946 XOR3X2 $T=1346400 1289680 0 0 $X=1346398 $Y=1289278
X1941 10329 10266 10238 1 3 8656 XOR3X2 $T=2030160 1188880 0 180 $X=2018280 $Y=1183440
X1942 10260 10297 10316 1 3 8627 XOR3X2 $T=2021580 1209040 0 0 $X=2021578 $Y=1208638
X1943 10502 10480 10476 1 3 8628 XOR3X2 $T=2062500 1269520 0 180 $X=2050620 $Y=1264080
X1944 10580 10572 10392 1 3 8173 XOR3X2 $T=2080320 1340080 1 180 $X=2068440 $Y=1339678
X1945 10609 562 10558 1 3 8168 XOR3X2 $T=2081640 1309840 1 180 $X=2069760 $Y=1309438
X1946 14256 691 14110 1 3 14106 XOR3X2 $T=2600400 1350160 0 180 $X=2588520 $Y=1344720
X1947 14127 693 692 1 3 14230 XOR3X2 $T=2593140 1400560 0 0 $X=2593138 $Y=1400158
X1948 1549 1664 3 1744 1 1808 AOI21XL $T=709500 1259440 0 0 $X=709498 $Y=1259038
X1949 1749 1807 3 1805 1 1778 AOI21XL $T=713460 1350160 1 180 $X=710820 $Y=1349758
X1950 1887 1807 3 1881 1 1611 AOI21XL $T=725340 1380400 0 180 $X=722700 $Y=1374960
X1951 2271 2270 3 2255 1 2207 AOI21XL $T=777480 1198960 0 180 $X=774840 $Y=1193520
X1952 2316 2270 3 2323 1 2349 AOI21XL $T=784080 1198960 1 0 $X=784078 $Y=1193520
X1953 5264 5262 3 253 1 5402 AOI21XL $T=1257300 1168720 1 0 $X=1257298 $Y=1163280
X1954 5459 5526 3 5542 1 5669 AOI21XL $T=1287660 1198960 1 0 $X=1287658 $Y=1193520
X1955 9381 9323 3 9353 1 9361 AOI21XL $T=1886280 1390480 1 180 $X=1883640 $Y=1390078
X1956 12746 12598 3 12723 1 12779 AOI21XL $T=2405700 1219120 0 0 $X=2405698 $Y=1218718
X1957 12835 637 3 12868 1 12895 AOI21XL $T=2424840 1158640 1 0 $X=2424838 $Y=1153200
X1958 13092 13183 3 13185 1 13189 AOI21XL $T=2472360 1400560 1 0 $X=2472358 $Y=1395120
X1959 654 13183 3 659 1 13428 AOI21XL $T=2502060 1420720 0 0 $X=2502058 $Y=1420318
X1960 13552 13183 3 13516 1 13520 AOI21XL $T=2517900 1410640 1 180 $X=2515260 $Y=1410238
X1961 13950 13902 3 13885 1 13906 AOI21XL $T=2564760 1158640 0 180 $X=2562120 $Y=1153200
X1962 14012 13942 3 14021 1 14033 AOI21XL $T=2575320 1269520 0 0 $X=2575318 $Y=1269118
X1963 696 14010 3 695 1 14334 AOI21XL $T=2618220 1410640 0 0 $X=2618218 $Y=1410238
X1964 1508 66 55 1 1599 3 OAI2BB1X1 $T=677820 1319920 1 0 $X=677818 $Y=1314480
X1965 1848 1752 1841 1 1805 3 OAI2BB1X1 $T=720060 1350160 1 180 $X=716760 $Y=1349758
X1966 3708 3586 3712 1 160 3 OAI2BB1X1 $T=1007160 1350160 0 0 $X=1007158 $Y=1349758
X1967 212 4434 4674 1 4614 3 OAI2BB1X1 $T=1166220 1420720 0 180 $X=1162920 $Y=1415280
X1968 192 4778 208 1 4849 3 OAI2BB1X1 $T=1191300 1138480 0 0 $X=1191298 $Y=1138078
X1969 4947 4953 4955 1 239 3 OAI2BB1X1 $T=1203180 1198960 0 0 $X=1203178 $Y=1198558
X1970 4857 4851 4987 1 5062 3 OAI2BB1X1 $T=1205820 1370320 1 0 $X=1205818 $Y=1364880
X1971 5109 5072 249 1 5135 3 OAI2BB1X1 $T=1224960 1289680 1 0 $X=1224958 $Y=1284240
X1972 5063 4954 5102 1 5220 3 OAI2BB1X1 $T=1229580 1188880 0 0 $X=1229578 $Y=1188478
X1973 5373 5375 5354 1 5351 3 OAI2BB1X1 $T=1255320 1229200 0 180 $X=1252020 $Y=1223760
X1974 5303 5226 5346 1 5487 3 OAI2BB1X1 $T=1257960 1198960 1 0 $X=1257958 $Y=1193520
X1975 5221 5356 5375 1 5435 3 OAI2BB1X1 $T=1260600 1239280 1 0 $X=1260598 $Y=1233840
X1976 5488 5553 5675 1 5716 3 OAI2BB1X1 $T=1309440 1158640 1 0 $X=1309438 $Y=1153200
X1977 6128 6088 6007 1 6260 3 OAI2BB1X1 $T=1387980 1330000 1 0 $X=1387978 $Y=1324560
X1978 6432 6309 6281 1 6406 3 OAI2BB1X1 $T=1434180 1229200 1 180 $X=1430880 $Y=1228798
X1979 6733 6796 6753 1 6826 3 OAI2BB1X1 $T=1488300 1289680 0 0 $X=1488298 $Y=1289278
X1980 8264 8245 8243 1 8363 3 OAI2BB1X1 $T=1707420 1309840 0 0 $X=1707418 $Y=1309438
X1981 524 9951 9792 1 9958 3 OAI2BB1X1 $T=1972080 1319920 1 0 $X=1972078 $Y=1314480
X1982 12402 626 12326 1 12327 3 OAI2BB1X1 $T=2360160 1410640 0 180 $X=2356860 $Y=1405200
X1983 12622 12395 12292 1 12773 3 OAI2BB1X1 $T=2400420 1209040 1 0 $X=2400418 $Y=1203600
X1984 12803 12572 12779 1 12905 3 OAI2BB1X1 $T=2423520 1219120 0 0 $X=2423518 $Y=1218718
X1985 13465 13339 13424 1 13432 3 OAI2BB1X1 $T=2508660 1188880 1 180 $X=2505360 $Y=1188478
X1986 1574 1 1576 3 1568 NAND2BXL $T=681780 1209040 1 0 $X=681778 $Y=1203600
X1987 2142 1 2145 3 1777 NAND2BXL $T=760320 1330000 1 180 $X=757680 $Y=1329598
X1988 2281 1 2285 3 2158 NAND2BXL $T=784080 1279600 1 180 $X=781440 $Y=1279198
X1989 2321 1 2346 3 2136 NAND2BXL $T=789360 1279600 0 180 $X=786720 $Y=1274160
X1990 3475 1 3465 3 3215 NAND2BXL $T=972180 1289680 1 180 $X=969540 $Y=1289278
X1991 3671 1 3615 3 3500 NAND2BXL $T=999900 1168720 1 180 $X=997260 $Y=1168318
X1992 3812 1 3836 3 3777 NAND2BXL $T=1029600 1330000 1 180 $X=1026960 $Y=1329598
X1993 177 1 206 3 4720 NAND2BXL $T=1181400 1380400 0 0 $X=1181398 $Y=1379998
X1994 196 1 252 3 5177 NAND2BXL $T=1236180 1410640 1 180 $X=1233540 $Y=1410238
X1995 6339 1 6379 3 6478 NAND2BXL $T=1424940 1410640 1 0 $X=1424938 $Y=1405200
X1996 7324 1 7286 3 7395 NAND2BXL $T=1576080 1340080 1 0 $X=1576078 $Y=1334640
X1997 7598 1 7625 3 7718 NAND2BXL $T=1618320 1249360 0 0 $X=1618318 $Y=1248958
X1998 11875 1 11853 3 11762 NAND2BXL $T=2280300 1410640 1 180 $X=2277660 $Y=1410238
X1999 11960 1 12040 3 12280 NAND2BXL $T=2337720 1299760 0 0 $X=2337718 $Y=1299358
X2000 12246 1 12185 3 12501 NAND2BXL $T=2346960 1269520 0 0 $X=2346958 $Y=1269118
X2001 653 1 652 3 13181 NAND2BXL $T=2488200 1390480 0 180 $X=2485560 $Y=1385040
X2002 4143 4095 4062 3922 3 1 3875 ADDFHX1 $T=1072500 1229200 1 180 $X=1057320 $Y=1228798
X2003 4205 4157 4125 3906 3 1 3951 ADDFHX1 $T=1083060 1340080 1 180 $X=1067880 $Y=1339678
X2004 4360 4301 4264 4209 3 1 4098 ADDFHX1 $T=1108140 1299760 0 180 $X=1092960 $Y=1294320
X2005 5946 299 6046 6045 3 1 6039 ADDFHX1 $T=1387320 1289680 1 180 $X=1372140 $Y=1289278
X2006 266 6127 6157 6160 3 1 6277 ADDFHX1 $T=1380060 1178800 1 0 $X=1380058 $Y=1173360
X2007 10529 549 10701 10702 3 1 10633 ADDFHX1 $T=2085600 1370320 1 0 $X=2085598 $Y=1364880
X2008 558 543 562 10946 3 1 11093 ADDFHX1 $T=2125860 1279600 0 0 $X=2125858 $Y=1279198
X2009 573 10172 10701 11147 3 1 11121 ADDFHX1 $T=2153580 1370320 0 0 $X=2153578 $Y=1369918
X2010 555 551 10520 11178 3 1 11486 ADDFHX1 $T=2162160 1259440 0 0 $X=2162158 $Y=1259038
X2011 605 609 570 11614 3 1 11625 ADDFHX1 $T=2230140 1168720 0 0 $X=2230138 $Y=1168318
X2012 11479 11732 11792 11805 3 1 11811 ADDFHX1 $T=2256540 1239280 0 0 $X=2256538 $Y=1238878
X2013 522 11598 11286 11810 3 1 11822 ADDFHX1 $T=2257860 1229200 1 0 $X=2257858 $Y=1223760
X2014 11814 11752 11804 11905 3 1 11908 ADDFHX1 $T=2273700 1148560 0 0 $X=2273698 $Y=1148158
X2015 4057 1 4030 3 4061 3921 NAND3X1 $T=1054680 1178800 0 180 $X=1052040 $Y=1173360
X2016 4152 1 4156 3 4177 4031 NAND3X1 $T=1074480 1269520 1 0 $X=1074478 $Y=1264080
X2017 4265 1 4262 3 4267 4215 NAND3X1 $T=1092300 1420720 0 180 $X=1089660 $Y=1415280
X2018 5839 1 5842 3 5832 5945 NAND3X1 $T=1345080 1249360 1 0 $X=1345078 $Y=1243920
X2019 7950 1 7953 3 7928 8013 NAND3X1 $T=1657260 1259440 0 0 $X=1657258 $Y=1259038
X2020 8164 1 8126 3 8241 8167 NAND3X1 $T=1698180 1239280 1 0 $X=1698178 $Y=1233840
X2021 8415 1 8362 3 8402 8430 NAND3X1 $T=1733160 1239280 1 0 $X=1733158 $Y=1233840
X2022 8401 1 8452 3 8144 8394 NAND3X1 $T=1737120 1168720 0 0 $X=1737118 $Y=1168318
X2023 9573 1 9570 3 9565 9563 NAND3X1 $T=1915320 1188880 1 180 $X=1912680 $Y=1188478
X2024 100 101 95 2487 1 3 2469 CMPR32X1 $T=818400 1410640 0 180 $X=804540 $Y=1405200
X2025 110 106 104 2522 1 3 2516 CMPR32X1 $T=827640 1360240 0 180 $X=813780 $Y=1354800
X2026 110 111 108 2489 1 3 2339 CMPR32X1 $T=845460 1420720 0 180 $X=831600 $Y=1415280
X2027 4214 4144 4098 4027 3 1 3957 ADDFHX2 $T=1085040 1299760 1 180 $X=1062600 $Y=1299358
X2028 4479 4484 4392 4450 3 1 4141 ADDFHX2 $T=1148400 1279600 1 180 $X=1125960 $Y=1279198
X2029 4511 4450 4457 3902 3 1 3903 ADDFHX2 $T=1149060 1259440 0 180 $X=1126620 $Y=1254000
X2030 5923 288 296 6036 3 1 6105 ADDFHX2 $T=1353000 1350160 0 0 $X=1352998 $Y=1349758
X2031 6257 5945 6045 6098 3 1 6087 ADDFHX2 $T=1403820 1269520 1 180 $X=1381380 $Y=1269118
X2032 268 6164 305 306 3 1 6335 ADDFHX2 $T=1389300 1158640 0 0 $X=1389298 $Y=1158238
X2033 6135 6191 6098 6309 3 1 6378 ADDFHX2 $T=1389960 1259440 0 0 $X=1389958 $Y=1259038
X2034 10529 11254 10302 11286 3 1 11479 ADDFHX2 $T=2176020 1229200 0 0 $X=2176018 $Y=1228798
X2035 11093 11283 11362 11387 3 1 11512 ADDFHX2 $T=2185260 1279600 0 0 $X=2185258 $Y=1279198
X2036 11486 11148 11606 11615 3 1 11553 ADDFHX2 $T=2222880 1289680 1 0 $X=2222878 $Y=1284240
X2037 610 11538 11625 11639 3 1 11698 ADDFHX2 $T=2226840 1188880 0 0 $X=2226838 $Y=1188478
X2038 11708 11787 11822 11827 3 1 12159 ADDFHX2 $T=2254560 1249360 0 0 $X=2254558 $Y=1248958
X2039 554 10676 558 10553 10558 1 3 ADDFHX4 $T=2108700 1279600 0 180 $X=2085600 $Y=1274160
X2040 58 55 1 3 1511 OR2X1 $T=663300 1269520 0 0 $X=663298 $Y=1269118
X2041 58 3 1602 1 CLKINVX3 $T=671880 1249360 0 0 $X=671878 $Y=1248958
X2042 118 3 3184 1 CLKINVX3 $T=920040 1400560 0 0 $X=920038 $Y=1400158
X2043 3371 3 3296 1 CLKINVX3 $T=953700 1259440 1 180 $X=951720 $Y=1259038
X2044 3437 3 3378 1 CLKINVX3 $T=960960 1299760 1 180 $X=958980 $Y=1299358
X2045 3416 3 3358 1 CLKINVX3 $T=967560 1299760 0 0 $X=967558 $Y=1299358
X2046 3816 3 3802 1 CLKINVX3 $T=1021680 1370320 1 180 $X=1019700 $Y=1369918
X2047 194 3 224 1 CLKINVX3 $T=1176120 1309840 1 180 $X=1174140 $Y=1309438
X2048 180 3 229 1 CLKINVX3 $T=1182060 1279600 0 0 $X=1182058 $Y=1279198
X2049 230 3 232 1 CLKINVX3 $T=1201860 1279600 0 180 $X=1199880 $Y=1274160
X2050 5498 3 6006 1 CLKINVX3 $T=1312740 1229200 1 0 $X=1312738 $Y=1223760
X2051 311 3 316 1 CLKINVX3 $T=1443420 1138480 0 0 $X=1443418 $Y=1138078
X2052 6946 3 6947 1 CLKINVX3 $T=1508760 1178800 0 0 $X=1508758 $Y=1178398
X2053 328 3 6998 1 CLKINVX3 $T=1511400 1289680 1 0 $X=1511398 $Y=1284240
X2054 7027 3 7031 1 CLKINVX3 $T=1524600 1239280 0 0 $X=1524598 $Y=1238878
X2055 336 3 326 1 CLKINVX3 $T=1547040 1430800 1 0 $X=1547038 $Y=1425360
X2056 7287 3 7478 1 CLKINVX3 $T=1568820 1198960 1 0 $X=1568818 $Y=1193520
X2057 357 3 7801 1 CLKINVX3 $T=1642080 1430800 1 0 $X=1642078 $Y=1425360
X2058 8117 3 8162 1 CLKINVX3 $T=1688940 1209040 0 0 $X=1688938 $Y=1208638
X2059 8187 3 8250 1 CLKINVX3 $T=1699500 1178800 0 0 $X=1699498 $Y=1178398
X2060 8782 3 430 1 CLKINVX3 $T=1793220 1148560 0 0 $X=1793218 $Y=1148158
X2061 8861 3 8864 1 CLKINVX3 $T=1801800 1340080 0 0 $X=1801798 $Y=1339678
X2062 8916 3 8954 1 CLKINVX3 $T=1824900 1350160 1 0 $X=1824898 $Y=1344720
X2063 9923 3 9854 1 CLKINVX3 $T=1968120 1249360 0 180 $X=1966140 $Y=1243920
X2064 9978 3 9897 1 CLKINVX3 $T=1978680 1239280 0 180 $X=1976700 $Y=1233840
X2065 10051 3 10141 1 CLKINVX3 $T=1997820 1269520 1 0 $X=1997818 $Y=1264080
X2066 10036 3 10143 1 CLKINVX3 $T=2008380 1269520 1 0 $X=2008378 $Y=1264080
X2067 10261 3 10207 1 CLKINVX3 $T=2022240 1309840 0 0 $X=2022238 $Y=1309438
X2068 566 3 556 1 CLKINVX3 $T=2079000 1370320 1 0 $X=2078998 $Y=1364880
X2069 11092 3 601 1 CLKINVX3 $T=2178660 1420720 0 0 $X=2178658 $Y=1420318
X2070 11451 3 11709 1 CLKINVX3 $T=2251260 1340080 0 0 $X=2251258 $Y=1339678
X2071 611 3 11734 1 CLKINVX3 $T=2263140 1390480 0 0 $X=2263138 $Y=1390078
X2072 12436 3 12598 1 CLKINVX3 $T=2379960 1239280 1 0 $X=2379958 $Y=1233840
X2073 12540 3 12632 1 CLKINVX3 $T=2387220 1370320 1 0 $X=2387218 $Y=1364880
X2074 13155 3 13159 1 CLKINVX3 $T=2465760 1269520 0 0 $X=2465758 $Y=1269118
X2075 13512 3 13508 1 CLKINVX3 $T=2514600 1289680 1 180 $X=2512620 $Y=1289278
X2076 13609 3 13514 1 CLKINVX3 $T=2525820 1239280 0 180 $X=2523840 $Y=1233840
X2077 13419 3 13312 1 CLKINVX3 $T=2530440 1229200 0 180 $X=2528460 $Y=1223760
X2078 13508 3 13698 1 CLKINVX3 $T=2533740 1279600 0 0 $X=2533738 $Y=1279198
X2079 1603 1655 3 1 1751 AND2X1 $T=691020 1209040 0 0 $X=691018 $Y=1208638
X2080 1807 1782 3 1 1672 AND2X1 $T=710820 1360240 0 180 $X=708180 $Y=1354800
X2081 3137 3197 3 1 3110 AND2X1 $T=933240 1158640 1 180 $X=930600 $Y=1158238
X2082 5922 5925 3 1 292 AND2X1 $T=1353660 1360240 0 0 $X=1353658 $Y=1359838
X2083 6737 6752 3 1 6870 AND2X1 $T=1479720 1158640 0 0 $X=1479718 $Y=1158238
X2084 11128 11094 3 1 599 AND2X1 $T=2167440 1430800 0 180 $X=2164800 $Y=1425360
X2085 12279 12424 3 1 12472 AND2X1 $T=2362140 1239280 0 0 $X=2362138 $Y=1238878
X2086 13610 13605 3 1 13650 AND2X1 $T=2535060 1299760 0 180 $X=2532420 $Y=1294320
X2087 13814 13813 3 1 13551 AND2X1 $T=2549580 1309840 0 180 $X=2546940 $Y=1304400
X2088 13816 13870 3 1 13805 AND2X1 $T=2552220 1410640 0 180 $X=2549580 $Y=1405200
X2089 13934 13927 3 1 13907 AND2X1 $T=2562780 1239280 1 180 $X=2560140 $Y=1238878
X2090 696 697 3 1 14336 AND2X1 $T=2607000 1420720 0 0 $X=2606998 $Y=1420318
X2091 1943 76 1954 3 1986 1 AOI2BB1X4 $T=731940 1350160 1 0 $X=731938 $Y=1344720
X2092 9721 9668 9766 3 9792 1 AOI2BB1X4 $T=1941060 1340080 0 0 $X=1941058 $Y=1339678
X2093 2305 2279 3 2330 2341 2353 1 AOI22X1 $T=784740 1219120 1 0 $X=784738 $Y=1213680
X2094 462 461 3 424 441 9043 1 AOI22X1 $T=1838760 1299760 1 180 $X=1835460 $Y=1299358
X2095 471 462 3 441 431 8975 1 AOI22X1 $T=1839420 1319920 0 180 $X=1836120 $Y=1314480
X2096 462 463 3 410 441 9062 1 AOI22X1 $T=1844700 1350160 0 180 $X=1841400 $Y=1344720
X2097 462 464 3 422 441 9038 1 AOI22X1 $T=1846020 1340080 1 180 $X=1842720 $Y=1339678
X2098 462 466 3 423 441 9068 1 AOI22X1 $T=1847340 1330000 0 180 $X=1844040 $Y=1324560
X2099 469 462 3 9328 441 9236 1 AOI22X1 $T=1884300 1269520 0 180 $X=1881000 $Y=1264080
X2100 472 462 3 9347 441 9297 1 AOI22X1 $T=1886940 1259440 0 180 $X=1883640 $Y=1254000
X2101 477 462 3 9386 441 9286 1 AOI22X1 $T=1892220 1239280 1 180 $X=1888920 $Y=1238878
X2102 494 462 3 9504 441 9405 1 AOI22X1 $T=1902120 1209040 0 180 $X=1898820 $Y=1203600
X2103 503 462 3 9443 441 9646 1 AOI22X1 $T=1928520 1148560 1 180 $X=1925220 $Y=1148158
X2104 507 462 3 9506 441 9723 1 AOI22X1 $T=1947000 1178800 0 180 $X=1943700 $Y=1173360
X2105 512 462 3 9508 441 9796 1 AOI22X1 $T=1950300 1209040 0 180 $X=1947000 $Y=1203600
X2106 10476 10480 3 10502 10501 10331 1 AOI22X1 $T=2061840 1259440 1 180 $X=2058540 $Y=1259038
X2107 10893 10889 3 10868 10890 10945 1 AOI22X1 $T=2131800 1410640 0 0 $X=2131798 $Y=1410238
X2108 14139 695 3 693 692 14226 1 AOI22X1 $T=2605680 1410640 1 180 $X=2602380 $Y=1410238
X2109 2380 2403 2313 2353 1 3 2255 OAI2BB2X1 $T=799260 1198960 0 180 $X=794640 $Y=1193520
X2110 182 4954 4947 177 1 3 4890 OAI2BB2X1 $T=1204500 1178800 0 180 $X=1199880 $Y=1173360
X2111 10299 10302 10298 10331 1 3 10325 OAI2BB2X1 $T=2038740 1239280 0 180 $X=2034120 $Y=1233840
X2112 10266 10238 10330 10356 1 3 10377 OAI2BB2X1 $T=2036760 1188880 1 0 $X=2036758 $Y=1183440
X2113 10531 10520 10530 10527 1 3 10502 OAI2BB2X1 $T=2067780 1279600 0 180 $X=2063160 $Y=1274160
X2114 562 10558 10607 10648 1 3 10632 OAI2BB2X1 $T=2090880 1330000 0 180 $X=2086260 $Y=1324560
X2115 104 87 95 2485 1 3 2514 ADDFXL $T=824340 1239280 0 180 $X=810480 $Y=1233840
X2116 97 87 1 3 2544 XNOR2XL $T=811140 1370320 1 0 $X=811138 $Y=1364880
X2117 110 108 1 3 2523 XNOR2XL $T=830940 1330000 1 180 $X=825660 $Y=1329598
X2118 5227 4990 1 3 5277 XNOR2XL $T=1238820 1279600 1 0 $X=1238818 $Y=1274160
X2119 5234 5277 1 3 5348 XNOR2XL $T=1246740 1279600 1 0 $X=1246738 $Y=1274160
X2120 188 210 1 3 5781 XNOR2XL $T=1327920 1330000 1 0 $X=1327918 $Y=1324560
X2121 2619 2171 2635 3 1 OR2X4 $T=834240 1188880 1 0 $X=834238 $Y=1183440
X2122 275 274 5587 3 1 OR2X4 $T=1299540 1360240 1 180 $X=1295580 $Y=1359838
X2123 3423 315 6572 3 1 OR2X4 $T=1451340 1360240 1 0 $X=1451338 $Y=1354800
X2124 6629 5994 6702 3 1 OR2X4 $T=1471140 1168720 0 0 $X=1471138 $Y=1168318
X2125 3359 321 6759 3 1 OR2X4 $T=1480380 1340080 1 0 $X=1480378 $Y=1334640
X2126 7000 3013 6978 3 1 OR2X4 $T=1518000 1219120 1 180 $X=1514040 $Y=1218718
X2127 7005 3355 6979 3 1 OR2X4 $T=1518000 1249360 0 180 $X=1514040 $Y=1243920
X2128 7095 6839 7103 3 1 OR2X4 $T=1534500 1350160 0 0 $X=1534498 $Y=1349758
X2129 7162 6725 7055 3 1 OR2X4 $T=1543080 1400560 0 0 $X=1543078 $Y=1400158
X2130 6922 7389 7392 3 1 OR2X4 $T=1574100 1299760 0 0 $X=1574098 $Y=1299358
X2131 7288 7760 7764 3 1 OR2X4 $T=1632180 1229200 1 0 $X=1632178 $Y=1223760
X2132 7655 7806 7837 3 1 OR2X4 $T=1642740 1198960 0 0 $X=1642738 $Y=1198558
X2133 447 448 8894 3 1 OR2X4 $T=1807080 1340080 0 0 $X=1807078 $Y=1339678
X2134 486 485 9381 3 1 OR2X4 $T=1894860 1390480 1 180 $X=1890900 $Y=1390078
X2135 500 499 9665 3 1 OR2X4 $T=1931160 1350160 0 180 $X=1927200 $Y=1344720
X2136 470 9692 9696 3 1 OR2X4 $T=1931160 1390480 0 0 $X=1931158 $Y=1390078
X2137 511 521 9903 3 1 OR2X4 $T=1964160 1360240 1 0 $X=1964158 $Y=1354800
X2138 619 12132 11928 3 1 OR2X4 $T=2321220 1390480 0 180 $X=2317260 $Y=1385040
X2139 646 13129 12999 3 1 OR2X4 $T=2465100 1330000 1 180 $X=2461140 $Y=1329598
X2140 2868 2789 2765 1 3 114 OAI2BB1X4 $T=859980 1178800 0 180 $X=853380 $Y=1173360
X2141 2916 2868 1 3 INVX8 $T=881100 1229200 1 180 $X=877140 $Y=1228798
X2142 3353 117 1 3 INVX8 $T=924660 1219120 0 180 $X=920700 $Y=1213680
X2143 10236 10076 1 3 INVX8 $T=2016960 1279600 0 180 $X=2013000 $Y=1274160
X2144 572 573 1 3 INVX8 $T=2093520 1380400 0 180 $X=2089560 $Y=1374960
X2145 11360 609 1 3 INVX8 $T=2212320 1209040 1 0 $X=2212318 $Y=1203600
X2146 13458 13222 1 3 INVX8 $T=2505360 1209040 1 0 $X=2505358 $Y=1203600
X2147 2874 2764 2872 2944 3 1 MX2X4 $T=882420 1178800 1 0 $X=882418 $Y=1173360
X2148 10144 532 10148 10172 3 1 MX2X4 $T=2000460 1420720 0 0 $X=2000458 $Y=1420318
X2149 2868 2953 2953 1 2868 3013 3 OAI2BB2X4 $T=889020 1219120 0 0 $X=889018 $Y=1218718
X2150 2898 2948 2986 1 3 NAND2BX2 $T=894960 1309840 0 0 $X=894958 $Y=1309438
X2151 2841 2946 3108 1 3 NAND2BX2 $T=900900 1269520 0 0 $X=900898 $Y=1269118
X2152 8860 8894 8942 1 3 NAND2BX2 $T=1815000 1360240 1 0 $X=1814998 $Y=1354800
X2153 3089 3065 3062 3061 3 1 OAI2BB1X2 $T=908820 1390480 1 180 $X=904200 $Y=1390078
X2154 174 171 4091 4051 3 1 OAI2BB1X2 $T=1065900 1430800 0 180 $X=1061280 $Y=1425360
X2155 13512 13605 13610 13548 3 1 OAI2BB1X2 $T=2523840 1299760 1 0 $X=2523838 $Y=1294320
X2156 13940 13698 13930 13911 3 1 OAI2BB1X2 $T=2564760 1279600 0 180 $X=2560140 $Y=1274160
X2157 134 136 3407 1 3 132 AND3X1 $T=963600 1178800 0 180 $X=960300 $Y=1173360
X2158 128 138 130 1 3 3407 AND3X2 $T=984720 1209040 1 180 $X=981420 $Y=1208638
X2159 336 7396 343 1 3 6440 AND3X2 $T=1578060 1420720 1 180 $X=1574760 $Y=1420318
X2160 434 7396 8750 1 3 436 AND3X2 $T=1788600 1410640 0 0 $X=1788598 $Y=1410238
X2161 142 1 3674 143 3 3670 NAND3BXL $T=1005180 1148560 0 180 $X=1001880 $Y=1143120
X2162 8043 1 350 372 3 374 NAND3BXL $T=1674420 1430800 1 0 $X=1674418 $Y=1425360
X2163 3615 3675 3595 1 3 NOR2BX2 $T=1005840 1178800 1 180 $X=1001880 $Y=1178398
X2164 6972 6976 6977 1 3 NOR2BX2 $T=1511400 1350160 1 0 $X=1511398 $Y=1344720
X2165 390 8271 8390 1 3 NOR2BX2 $T=1717980 1420720 1 0 $X=1717978 $Y=1415280
X2166 8120 8271 8379 1 3 NOR2BX2 $T=1725240 1390480 0 0 $X=1725238 $Y=1390078
X2167 14313 12493 14073 1 3 NOR2BX2 $T=2618880 1239280 0 0 $X=2618878 $Y=1238878
X2168 166 165 1 3 3534 XOR2XL $T=1021680 1410640 1 180 $X=1016400 $Y=1410238
X2169 5072 5241 1 3 5492 XOR2XL $T=1240800 1289680 0 0 $X=1240798 $Y=1289278
X2170 391 8397 1 3 8400 XOR2XL $T=1738440 1138480 1 180 $X=1733160 $Y=1138078
X2171 8491 8632 1 3 8618 XOR2XL $T=1767480 1289680 1 180 $X=1762200 $Y=1289278
X2172 431 9558 1 3 9507 XOR2XL $T=1911360 1279600 1 180 $X=1906080 $Y=1279198
X2173 3 4439 4144 4411 4455 1 NAND3X2 $T=1121340 1319920 0 0 $X=1121338 $Y=1319518
X2174 3 9708 9401 9712 9621 1 NAND3X2 $T=1937760 1289680 1 180 $X=1933140 $Y=1289278
X2175 3 9872 9591 9702 9740 1 NAND3X2 $T=1935120 1269520 0 0 $X=1935118 $Y=1269118
X2176 202 203 4434 4435 207 3 1 4464 SDFFRHQXL $T=1122000 1410640 0 0 $X=1121998 $Y=1410238
X2177 202 203 189 4524 207 3 1 4467 SDFFRHQXL $T=1147740 1410640 0 180 $X=1131240 $Y=1405200
X2178 202 203 235 233 207 3 1 4818 SDFFRHQXL $T=1206480 1410640 0 180 $X=1189980 $Y=1405200
X2179 202 203 177 238 207 3 1 4812 SDFFRHQXL $T=1211100 1430800 0 180 $X=1194600 $Y=1425360
X2180 202 203 179 4753 207 3 1 5523 SDFFRHQXL $T=1268520 1410640 1 0 $X=1268518 $Y=1405200
X2181 202 203 272 5188 207 3 1 5099 SDFFRHQXL $T=1289640 1410640 0 0 $X=1289638 $Y=1410238
X2182 202 203 5099 281 207 3 1 5612 SDFFRHQXL $T=1316040 1410640 0 180 $X=1299540 $Y=1405200
X2183 347 349 350 7620 354 3 1 7465 SDFFRHQXL $T=1603800 1420720 1 0 $X=1603798 $Y=1415280
X2184 347 349 7465 7627 354 3 1 7521 SDFFRHQXL $T=1605780 1400560 1 0 $X=1605778 $Y=1395120
X2185 347 349 7521 7648 354 3 1 7523 SDFFRHQXL $T=1609080 1360240 0 0 $X=1609078 $Y=1359838
X2186 347 349 7523 7654 354 3 1 7526 SDFFRHQXL $T=1609740 1350160 1 0 $X=1609738 $Y=1344720
X2187 347 349 7526 7786 354 3 1 7821 SDFFRHQXL $T=1633500 1340080 1 0 $X=1633498 $Y=1334640
X2188 347 349 7821 8007 354 3 1 368 SDFFRHQXL $T=1663200 1340080 1 0 $X=1663198 $Y=1334640
X2189 347 349 368 8041 354 3 1 7838 SDFFRHQXL $T=1680360 1319920 0 180 $X=1663860 $Y=1314480
X2190 347 349 7920 8013 354 3 1 7924 SDFFRHQXL $T=1666500 1279600 0 0 $X=1666498 $Y=1279198
X2191 347 349 7838 8015 354 3 1 7920 SDFFRHQXL $T=1666500 1299760 0 0 $X=1666498 $Y=1299358
X2192 347 349 7924 8167 354 3 1 8242 SDFFRHQXL $T=1692240 1259440 0 0 $X=1692238 $Y=1259038
X2193 347 349 8242 8430 354 3 1 8311 SDFFRHQXL $T=1738440 1259440 1 180 $X=1721940 $Y=1259038
X2194 347 349 8277 8342 354 3 1 8335 SDFFRHQXL $T=1722600 1219120 1 0 $X=1722598 $Y=1213680
X2195 347 349 8311 8361 354 3 1 8277 SDFFRHQXL $T=1722600 1239280 0 0 $X=1722598 $Y=1238878
X2196 454 453 422 8949 446 3 1 423 SDFFRHQXL $T=1822260 1430800 0 180 $X=1805760 $Y=1425360
X2197 347 453 461 9076 446 3 1 9230 SDFFRHQXL $T=1845360 1279600 0 0 $X=1845358 $Y=1279198
X2198 347 453 469 8984 446 3 1 9229 SDFFRHQXL $T=1846020 1269520 1 0 $X=1846018 $Y=1264080
X2199 347 453 472 9207 446 3 1 9111 SDFFRHQXL $T=1862520 1239280 0 180 $X=1846020 $Y=1233840
X2200 347 453 463 9209 446 3 1 422 SDFFRHQXL $T=1863180 1360240 1 180 $X=1846680 $Y=1359838
X2201 347 453 464 8977 446 3 1 9262 SDFFRHQXL $T=1849980 1309840 0 0 $X=1849978 $Y=1309438
X2202 347 453 431 9130 446 3 1 9244 SDFFRHQXL $T=1850640 1299760 0 0 $X=1850638 $Y=1299358
X2203 347 453 471 9058 446 3 1 9266 SDFFRHQXL $T=1851300 1340080 1 0 $X=1851298 $Y=1334640
X2204 347 453 477 9327 446 3 1 9205 SDFFRHQXL $T=1884300 1229200 1 180 $X=1867800 $Y=1228798
X2205 347 453 9347 9343 446 3 1 9269 SDFFRHQXL $T=1885620 1219120 1 180 $X=1869120 $Y=1218718
X2206 347 453 9328 9399 446 3 1 431 SDFFRHQXL $T=1895520 1309840 0 180 $X=1879020 $Y=1304400
X2207 347 453 466 9401 446 3 1 9328 SDFFRHQXL $T=1896180 1299760 0 180 $X=1879680 $Y=1294320
X2208 347 453 9386 9591 446 3 1 9347 SDFFRHQXL $T=1921260 1269520 1 180 $X=1904760 $Y=1269118
X2209 347 453 495 9404 446 3 1 497 SDFFRHQXL $T=1906080 1158640 1 0 $X=1906078 $Y=1153200
X2210 347 453 494 9563 446 3 1 9443 SDFFRHQXL $T=1907400 1168720 0 0 $X=1907398 $Y=1168318
X2211 347 453 9504 9617 446 3 1 9386 SDFFRHQXL $T=1924560 1239280 1 180 $X=1908060 $Y=1238878
X2212 347 453 9508 9634 446 3 1 9504 SDFFRHQXL $T=1927860 1229200 0 180 $X=1911360 $Y=1223760
X2213 347 453 9443 9728 446 3 1 9813 SDFFRHQXL $T=1933800 1168720 1 0 $X=1933798 $Y=1163280
X2214 347 453 507 9790 446 3 1 495 SDFFRHQXL $T=1950960 1158640 1 180 $X=1934460 $Y=1158238
X2215 347 453 503 9738 446 3 1 9850 SDFFRHQXL $T=1935780 1148560 0 0 $X=1935778 $Y=1148158
X2216 347 453 9506 9772 446 3 1 9508 SDFFRHQXL $T=1940400 1219120 0 0 $X=1940398 $Y=1218718
X2217 347 453 512 9763 446 3 1 9506 SDFFRHQXL $T=1956900 1209040 1 180 $X=1940400 $Y=1208638
X2218 4464 3 206 1 BUFX3 $T=1131240 1400560 0 180 $X=1128600 $Y=1395120
X2219 4467 3 4434 1 BUFX3 $T=1137840 1400560 1 0 $X=1137838 $Y=1395120
X2220 221 3 208 1 BUFX3 $T=1166220 1209040 1 0 $X=1166218 $Y=1203600
X2221 196 3 228 1 BUFX3 $T=1179420 1269520 1 0 $X=1179418 $Y=1264080
X2222 5431 3 5434 1 BUFX3 $T=1267200 1360240 1 0 $X=1267198 $Y=1354800
X2223 348 3 350 1 BUFX3 $T=1609080 1430800 1 0 $X=1609078 $Y=1425360
X2224 7527 3 379 1 BUFX3 $T=1690920 1188880 0 0 $X=1690918 $Y=1188478
X2225 7479 3 8149 1 BUFX3 $T=1691580 1219120 0 0 $X=1691578 $Y=1218718
X2226 8271 3 389 1 BUFX3 $T=1717980 1269520 0 180 $X=1715340 $Y=1264080
X2227 8618 3 425 1 BUFX3 $T=1762200 1309840 0 0 $X=1762198 $Y=1309438
X2228 8684 3 427 1 BUFX3 $T=1775400 1259440 1 0 $X=1775398 $Y=1254000
X2229 8271 3 462 1 BUFX3 $T=1824900 1269520 0 0 $X=1824898 $Y=1269118
X2230 9111 3 469 1 BUFX3 $T=1854600 1229200 0 0 $X=1854598 $Y=1228798
X2231 9205 3 472 1 BUFX3 $T=1857240 1219120 1 180 $X=1854600 $Y=1218718
X2232 9229 3 461 1 BUFX3 $T=1857240 1259440 0 180 $X=1854600 $Y=1254000
X2233 9262 3 471 1 BUFX3 $T=1861200 1319920 1 180 $X=1858560 $Y=1319518
X2234 9244 3 464 1 BUFX3 $T=1865160 1309840 1 0 $X=1865158 $Y=1304400
X2235 9230 3 466 1 BUFX3 $T=1867800 1279600 0 0 $X=1867798 $Y=1279198
X2236 9269 3 477 1 BUFX3 $T=1873080 1209040 0 0 $X=1873078 $Y=1208638
X2237 9266 3 463 1 BUFX3 $T=1884960 1340080 1 0 $X=1884958 $Y=1334640
X2238 449 3 9868 1 BUFX3 $T=1955580 1299760 0 0 $X=1955578 $Y=1299358
X2239 9813 3 512 1 BUFX3 $T=1956900 1168720 1 0 $X=1956898 $Y=1163280
X2240 9850 3 507 1 BUFX3 $T=1959540 1148560 0 0 $X=1959538 $Y=1148158
X2241 10521 3 560 1 BUFX3 $T=2063820 1370320 0 0 $X=2063818 $Y=1369918
X2242 10172 3 557 1 BUFX3 $T=2115960 1219120 0 180 $X=2113320 $Y=1213680
X2243 11707 3 12572 1 BUFX3 $T=2391840 1299760 1 0 $X=2391838 $Y=1294320
X2244 215 216 217 3 177 1 4538 4438 AOI221X1 $T=1147740 1420720 0 0 $X=1147738 $Y=1420318
X2245 4617 219 192 3 4615 184 1 4670 AOI32XL $T=1153680 1370320 1 0 $X=1153678 $Y=1364880
X2246 4307 222 4720 3 177 4725 1 4724 AOI32XL $T=1168860 1380400 0 0 $X=1168858 $Y=1379998
X2247 5103 246 189 3 242 187 1 5143 AOI32XL $T=1223640 1410640 0 0 $X=1223638 $Y=1410238
X2248 198 256 5177 3 196 255 1 5198 AOI32XL $T=1244100 1410640 1 180 $X=1239480 $Y=1410238
X2249 5944 5948 128 3 5849 138 1 6029 AOI32XL $T=1358280 1410640 1 0 $X=1358278 $Y=1405200
X2250 5998 6002 134 3 6028 136 1 6030 AOI32XL $T=1367520 1390480 0 0 $X=1367518 $Y=1390078
X2251 6190 5948 197 3 6123 179 1 6193 AOI32XL $T=1403160 1390480 0 180 $X=1398540 $Y=1385040
X2252 9204 9187 479 3 9188 470 1 9441 AOI32XL $T=1885620 1430800 1 0 $X=1885618 $Y=1425360
X2253 221 205 3 1 CLKINVX4 $T=1164900 1219120 0 0 $X=1164898 $Y=1218718
X2254 216 162 3 225 217 212 223 4726 1 AOI222X2 $T=1180740 1420720 1 180 $X=1171500 $Y=1420318
X2255 204 4807 1 4665 189 3 4811 OAI22X1 $T=1191300 1198960 0 180 $X=1187340 $Y=1193520
X2256 4807 4844 1 4665 208 3 4953 OAI22X1 $T=1193940 1198960 1 180 $X=1189980 $Y=1198558
X2257 231 3 209 4948 1 NOR2BXL $T=1194600 1340080 0 0 $X=1194598 $Y=1339678
X2258 244 3 180 5071 1 NOR2BXL $T=1226940 1350160 1 180 $X=1224300 $Y=1349758
X2259 4857 3 4722 4881 1 4959 NOR3BX1 $T=1195260 1370320 1 0 $X=1195258 $Y=1364880
X2260 236 3 234 4949 1 4948 4857 AOI211X1 $T=1203840 1350160 0 180 $X=1200540 $Y=1344720
X2261 5305 3 5281 5213 1 5243 5267 AOI211X1 $T=1248720 1400560 1 180 $X=1245420 $Y=1400158
X2262 4948 236 234 1 231 240 3 4989 OAI32X1 $T=1206480 1340080 0 0 $X=1206478 $Y=1339678
X2263 5071 245 224 1 244 229 3 4991 OAI32X1 $T=1220340 1360240 0 180 $X=1215720 $Y=1354800
X2264 5267 5222 5062 1 4959 5062 3 5197 OAI32X1 $T=1240140 1370320 1 180 $X=1235520 $Y=1369918
X2265 5374 260 247 1 259 230 3 5347 OAI32X1 $T=1257300 1390480 0 180 $X=1252680 $Y=1385040
X2266 5032 4986 1 3 5023 267 AOI2BB1X1 $T=1219020 1148560 1 0 $X=1219018 $Y=1143120
X2267 329 7092 1 3 7133 7266 AOI2BB1X1 $T=1539120 1380400 0 0 $X=1539118 $Y=1379998
X2268 7358 6998 1 3 7383 7376 AOI2BB1X1 $T=1572120 1239280 1 0 $X=1572118 $Y=1233840
X2269 653 647 1 3 13282 13308 AOI2BB1X1 $T=2487540 1410640 1 0 $X=2487538 $Y=1405200
X2270 216 248 3 212 5099 189 5110 217 1 AOI222X1 $T=1225620 1420720 1 180 $X=1220340 $Y=1420318
X2271 7454 7479 3 7527 7295 7465 7513 7503 1 AOI222X1 $T=1599180 1400560 1 180 $X=1593900 $Y=1400158
X2272 7552 7479 3 7527 7512 7521 7553 7503 1 AOI222X1 $T=1599840 1390480 0 180 $X=1594560 $Y=1385040
X2273 7550 7479 3 7527 7531 7526 7544 7503 1 AOI222X1 $T=1601160 1340080 1 180 $X=1595880 $Y=1339678
X2274 7532 7479 3 7527 7472 7523 7558 7503 1 AOI222X1 $T=1601160 1360240 1 180 $X=1595880 $Y=1359838
X2275 7841 7479 3 7527 7753 7821 7798 7802 1 AOI222X1 $T=1646040 1309840 1 180 $X=1640760 $Y=1309438
X2276 7829 7479 3 7527 7792 7838 8016 7802 1 AOI222X1 $T=1651980 1309840 1 0 $X=1651978 $Y=1304400
X2277 7925 7479 3 7527 7921 7802 7927 7920 1 AOI222X1 $T=1657260 1289680 0 180 $X=1651980 $Y=1284240
X2278 411 8375 3 8379 262 304 8591 8390 1 AOI222X1 $T=1740420 1410640 0 0 $X=1740418 $Y=1410238
X2279 218 5185 254 5108 1 3 MXI2X1 $T=1234200 1239280 1 0 $X=1234198 $Y=1233840
X2280 5376 5353 1 5236 3 5345 5350 OAI211X1 $T=1254000 1158640 0 180 $X=1250040 $Y=1153200
X2281 5354 4811 1 5356 3 5221 5382 OAI211X1 $T=1261920 1229200 1 180 $X=1257960 $Y=1228798
X2282 5487 5488 1 5553 3 5485 271 OAI211X1 $T=1288980 1148560 0 0 $X=1288978 $Y=1148158
X2283 5487 5488 1 5485 3 5553 277 OAI211X1 $T=1303500 1148560 1 180 $X=1299540 $Y=1148158
X2284 8247 8250 1 8249 3 8175 8342 OAI211X1 $T=1701480 1209040 1 0 $X=1701478 $Y=1203600
X2285 9897 9853 1 9867 3 9871 9772 OAI211X1 $T=1962840 1229200 1 180 $X=1958880 $Y=1228798
X2286 5276 257 5221 1 3 5411 XNOR3X2 $T=1252680 1249360 1 0 $X=1252678 $Y=1243920
X2287 5191 5548 5526 1 3 5588 XNOR3X2 $T=1283040 1219120 1 0 $X=1283038 $Y=1213680
X2288 5520 5220 5669 1 3 5673 XNOR3X2 $T=1298220 1188880 1 0 $X=1298218 $Y=1183440
X2289 10265 538 10322 1 3 8919 XNOR3X2 $T=2022900 1138480 0 0 $X=2022898 $Y=1138078
X2290 10331 10299 10302 1 3 8863 XNOR3X2 $T=2041380 1249360 0 180 $X=2029500 $Y=1243920
X2291 10527 10531 10520 1 3 8574 XNOR3X2 $T=2073060 1289680 1 180 $X=2061180 $Y=1289278
X2292 188 3 5377 191 261 5281 1 AOI22XL $T=1258620 1410640 0 180 $X=1255320 $Y=1405200
X2293 261 191 1 262 3 5377 AOI2BB1XL $T=1255980 1410640 0 0 $X=1255978 $Y=1410238
X2294 5353 5376 3 5402 1 5236 5433 AOI211X2 $T=1257960 1158640 1 0 $X=1257958 $Y=1153200
X2295 5375 5373 1 3 5382 5351 5526 OAI211X2 $T=1261920 1219120 0 0 $X=1261918 $Y=1218718
X2296 5220 5520 1 3 5459 5526 5582 OAI211X2 $T=1290960 1188880 1 180 $X=1284360 $Y=1188478
X2297 5605 5650 1 3 5582 5584 5553 OAI211X2 $T=1300200 1178800 0 180 $X=1293600 $Y=1173360
X2298 9853 9854 1 3 9757 9773 9617 OAI211X2 $T=1953600 1239280 1 180 $X=1947000 $Y=1238878
X2299 263 3 264 101 265 5431 1 NOR4BX1 $T=1263240 1360240 1 0 $X=1263238 $Y=1354800
X2300 5485 5487 5488 5489 3 1 269 AOI31X4 $T=1277100 1148560 0 0 $X=1277098 $Y=1148158
X2301 5523 223 1 3 BUFX4 $T=1285020 1410640 1 0 $X=1285018 $Y=1405200
X2302 5612 179 1 3 BUFX4 $T=1307460 1400560 1 0 $X=1307458 $Y=1395120
X2303 7922 364 1 3 BUFX4 $T=1654620 1390480 0 0 $X=1654618 $Y=1390078
X2304 433 8780 1 3 BUFX4 $T=1790580 1400560 0 0 $X=1790578 $Y=1400158
X2305 11254 608 1 3 BUFX4 $T=2212320 1138480 0 0 $X=2212318 $Y=1138078
X2306 5555 104 273 1 97 3 5586 OR4X2 $T=1291620 1340080 0 0 $X=1291618 $Y=1339678
X2307 9033 457 9036 1 458 3 8949 OR4X2 $T=1830180 1420720 0 0 $X=1830178 $Y=1420318
X2308 523 518 517 1 516 3 9722 OR4X2 $T=1961520 1430800 0 180 $X=1957560 $Y=1425360
X2309 5587 5434 1 3 5555 NAND2BX4 $T=1299540 1350160 0 180 $X=1294260 $Y=1344720
X2310 9069 9322 1 3 9317 NAND2BX4 $T=1879680 1380400 0 180 $X=1874400 $Y=1374960
X2311 10349 10295 1 3 10235 NAND2BX4 $T=2029500 1330000 1 180 $X=2024220 $Y=1329598
X2312 296 5973 284 5835 3 1 ADDHX4 $T=1372140 1279600 1 180 $X=1353660 $Y=1279198
X2313 6001 6002 200 3 6028 298 1 6040 AOI32X1 $T=1368180 1370320 0 0 $X=1368178 $Y=1369918
X2314 669 667 13816 3 672 670 1 13877 AOI32X1 $T=2546940 1420720 0 0 $X=2546938 $Y=1420318
X2315 297 5972 1 6089 6066 6100 6106 3 302 OAI33X1 $T=1380060 1420720 1 0 $X=1380058 $Y=1415280
X2316 5197 6365 1 6366 6343 6370 6371 3 309 OAI33X1 $T=1419660 1370320 0 0 $X=1419658 $Y=1369918
X2317 6106 6100 5999 3 1 6089 OR3XL $T=1384680 1410640 0 180 $X=1381380 $Y=1405200
X2318 6371 6370 6250 3 1 6366 OR3XL $T=1424940 1360240 1 180 $X=1421640 $Y=1359838
X2319 520 518 516 3 1 10177 OR3XL $T=2019600 1400560 0 180 $X=2016300 $Y=1395120
X2320 7283 7349 1 6998 7328 7348 3 OAI22XL $T=1568160 1239280 1 180 $X=1564200 $Y=1238878
X2321 7282 6998 338 1 7379 3 7388 OAI31X1 $T=1569480 1269520 0 0 $X=1569478 $Y=1269118
X2322 7396 7466 343 7479 1 3 AND3X4 $T=1587300 1420720 1 0 $X=1587298 $Y=1415280
X2323 433 7396 8750 435 1 3 AND3X4 $T=1786620 1400560 0 0 $X=1786618 $Y=1400158
X2324 3 7465 7521 7523 7526 7754 1 NOR4X1 $T=1637460 1390480 1 0 $X=1637458 $Y=1385040
X2325 3 7465 7521 7523 7526 7795 1 NOR4X1 $T=1641420 1380400 1 180 $X=1637460 $Y=1379998
X2326 3 7821 7838 7920 7924 7930 1 NOR4X1 $T=1655280 1370320 1 0 $X=1655278 $Y=1364880
X2327 3 7821 7838 7920 7924 7771 1 NOR4X1 $T=1665180 1370320 1 0 $X=1665178 $Y=1364880
X2328 3 8373 8303 392 391 8340 1 NOR4X1 $T=1721940 1340080 0 180 $X=1717980 $Y=1334640
X2329 3 8242 8311 8277 8335 8381 1 NOR4X1 $T=1728540 1309840 1 180 $X=1724580 $Y=1309438
X2330 3 8242 8311 8277 8335 8338 1 NOR4X1 $T=1725900 1319920 0 0 $X=1725898 $Y=1319518
X2331 3 8373 8303 392 391 8413 1 NOR4X1 $T=1731180 1330000 0 0 $X=1731178 $Y=1329598
X2332 3 9443 9504 9506 9508 9324 1 NOR4X1 $T=1898820 1219120 1 0 $X=1898818 $Y=1213680
X2333 3 9443 9504 9506 9508 9444 1 NOR4X1 $T=1898820 1229200 1 0 $X=1898818 $Y=1223760
X2334 363 1 367 3 361 7989 NAND3XL $T=1669140 1400560 1 180 $X=1666500 $Y=1400158
X2335 362 370 3 367 363 1 373 8043 AOI221XL $T=1673760 1420720 1 0 $X=1673758 $Y=1415280
X2336 368 367 363 1 7951 3 OAI2BB1XL $T=1677720 1400560 1 180 $X=1674420 $Y=1400158
X2337 8244 8166 1 8188 8251 3 8247 8162 8361 OAI222X1 $T=1700160 1209040 0 0 $X=1700158 $Y=1208638
X2338 384 1 8271 3 CLKINVX8 $T=1704120 1430800 0 180 $X=1700160 $Y=1425360
X2339 8271 3 363 1 377 8265 NOR3X1 $T=1707420 1410640 1 180 $X=1704780 $Y=1410238
X2340 8375 402 8379 272 8390 7526 393 1 3 AOI222X4 $T=1729860 1410640 0 180 $X=1721940 $Y=1405200
X2341 8375 394 8379 258 8390 7465 417 1 3 AOI222X4 $T=1722600 1400560 0 0 $X=1722598 $Y=1400158
X2342 8379 231 8375 399 8311 8390 8414 1 3 AOI222X4 $T=1723920 1340080 0 0 $X=1723918 $Y=1339678
X2343 8375 395 8379 206 8390 7838 407 1 3 AOI222X4 $T=1723920 1370320 0 0 $X=1723918 $Y=1369918
X2344 8375 396 8379 223 7821 8390 405 1 3 AOI222X4 $T=1723920 1380400 0 0 $X=1723918 $Y=1379998
X2345 8379 245 8375 400 8277 8390 8417 1 3 AOI222X4 $T=1724580 1350160 1 0 $X=1724578 $Y=1344720
X2346 8379 213 8375 403 7924 8390 406 1 3 AOI222X4 $T=1726560 1370320 1 0 $X=1726558 $Y=1364880
X2347 8375 401 8379 404 303 8390 8433 1 3 AOI222X4 $T=1727220 1420720 1 0 $X=1727218 $Y=1415280
X2348 8379 304 8375 410 8373 8390 8679 1 3 AOI222X4 $T=1737120 1360240 1 0 $X=1737118 $Y=1354800
X2349 8375 408 8379 5099 8390 7523 415 1 3 AOI222X4 $T=1737120 1410640 1 0 $X=1737118 $Y=1405200
X2350 8379 236 8375 412 8242 8390 8498 1 3 AOI222X4 $T=1739760 1340080 0 0 $X=1739758 $Y=1339678
X2351 8379 4434 8375 413 7920 8390 416 1 3 AOI222X4 $T=1739760 1370320 0 0 $X=1739758 $Y=1369918
X2352 8379 244 8375 414 8335 8390 8575 1 3 AOI222X4 $T=1740420 1350160 1 0 $X=1740418 $Y=1344720
X2353 8375 419 8379 260 314 8390 8625 1 3 AOI222X4 $T=1749000 1380400 0 0 $X=1748998 $Y=1379998
X2354 8375 421 8379 252 8390 7521 418 1 3 AOI222X4 $T=1756920 1390480 1 180 $X=1749000 $Y=1390078
X2355 8375 420 8379 259 325 8390 8649 1 3 AOI222X4 $T=1753620 1410640 1 0 $X=1753618 $Y=1405200
X2356 8379 314 8375 423 392 8390 8596 1 3 AOI222X4 $T=1754280 1350160 1 0 $X=1754278 $Y=1344720
X2357 325 8379 422 8375 8390 391 8619 1 3 AOI222X4 $T=1754280 1370320 0 0 $X=1754278 $Y=1369918
X2358 8379 303 8375 424 8303 8390 8620 1 3 AOI222X4 $T=1754940 1340080 1 0 $X=1754938 $Y=1334640
X2359 347 349 8335 8394 354 8451 1 3 8373 SDFFRXL $T=1722600 1178800 1 0 $X=1722598 $Y=1173360
X2360 347 349 8451 8148 354 397 1 3 8303 SDFFRXL $T=1741740 1158640 1 180 $X=1723260 $Y=1158238
X2361 433 356 3 1 449 NOR2BX4 $T=1797180 1390480 1 0 $X=1797178 $Y=1385040
X2362 9122 1 467 9103 9065 9189 3 NOR4X2 $T=1844040 1410640 1 0 $X=1844038 $Y=1405200
X2363 9386 3 9347 9328 431 9326 1 NOR4XL $T=1892220 1269520 1 180 $X=1888260 $Y=1269118
X2364 9386 3 9347 9328 431 9437 1 NOR4XL $T=1900140 1269520 0 180 $X=1896180 $Y=1264080
X2365 9722 504 502 501 1 9692 3 NAND4BBX2 $T=1937100 1430800 0 180 $X=1929840 $Y=1425360
X2366 9763 9756 9771 3 1 9739 NAND3BX2 $T=1945020 1198960 0 180 $X=1939740 $Y=1193520
X2367 9853 514 8780 1 510 3 9791 509 9790 OAI222XL $T=1954260 1148560 0 180 $X=1948980 $Y=1143120
X2368 521 511 1 3 9920 AND2X4 $T=1962840 1350160 0 0 $X=1962838 $Y=1349758
X2369 527 526 1 3 9959 AND2X4 $T=1986600 1360240 0 0 $X=1986598 $Y=1359838
X2370 13507 13504 1 3 13415 AND2X4 $T=2514600 1229200 0 180 $X=2511300 $Y=1223760
X2371 10177 523 533 1 3 10208 MX2X1 $T=2009700 1390480 1 0 $X=2009698 $Y=1385040
X2372 10208 543 1 3 INVX12 $T=2015640 1390480 1 0 $X=2015638 $Y=1385040
X2373 12038 3 1 7095 BUFX8 $T=2301420 1350160 1 180 $X=2295480 $Y=1349758
X2374 12271 12272 3 12159 11805 12273 1 AOI22X2 $T=2343000 1279600 0 180 $X=2337060 $Y=1274160
X2375 12876 7389 1 3 BUFX16 $T=2429460 1309840 1 0 $X=2429458 $Y=1304400
X2376 13419 657 13415 13312 1 3 MXI2X4 $T=2503380 1229200 0 180 $X=2494140 $Y=1223760
.ENDS
***************************************
.SUBCKT OAI211XL A1 A0 VSS C0 VDD B0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRHQX1 CK SE SI D RN VDD VSS Q
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ANTENNA VSS VDD A
** N=5 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRHQX2 CK SE SI D RN Q VSS VDD
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX12 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRHQX4 CK SI SE D RN VDD VSS Q
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB2XL A1N A0N B1 VDD B0 Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221X4 B1 B0 A0 A1 C0 Y VDD VSS
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222X4 B1 B0 A0 A1 C1 C0 Y VDD VSS
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221X1 B1 B0 A0 VSS A1 VDD C0 Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRX4 CK SE SI D RN QN Q VSS VDD
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4X1 D VSS C B A Y VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22X4 B0 VDD B1 A1 VSS A0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22X2 B1 VSS B0 A1 VDD A0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFXL A VSS VDD Y
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI31X2 A2 A1 A0 VDD B0 Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3X4 C VSS B A VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3BX1 AN VSS C B VDD Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22X4 B0 VSS B1 VDD A1 A0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX2 A VDD VSS Y
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3X4 A B C Y VSS VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR3X4 B C VDD VSS A Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX2 A VSS Y VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221X2 B1 B0 VSS A0 A1 C0 VDD Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX20 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4X4 A B C D VDD VSS Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI221X2 B0 B1 VDD A1 A0 VSS C0 Y
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MX2X2 B S0 A VDD VSS Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI211XL A1 A0 VDD C0 VSS B0 Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI2X2 S0 B Y A VSS VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_60 1 2 3 21 22 24 25 26 27 28 29 30 31 33 34 35 37 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 57 59 60 61 63 64 65
+ 66 67 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106
+ 107 108 109 110 111 112 114 115 117 118 119 120 122 123 124 125 126 128 129 130
+ 131 133 134 135 137 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153
+ 154 155 156 157 159 160 161 163 164 165 167 168 169 170 171 173 174 175 176 178
+ 179 180 181 182 183 184 185 186 188 189 190 191 192 193 194 195 196 197 198 199
+ 200 201 202 203 204 205 206 207 208 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 229 230 231 232 233 234 235 236 237 238 239 240 242
+ 243 244 245 247 248 249 250 251 252 254 255 256 257 258 259 260 261 262 263 264
+ 265 267 268 270 271 272 273 274 275 276 278 280 281 282 283 284 285 286 287 288
+ 289 290 291 292 293 295 296 298 300 301 302 303 304 305 307 308 309 311 313 314
+ 315 316 317 318 320 321 323 324 325 327 329 330 331 332 333 335 336 337 339 340
+ 341 342 344 346 347 348 349 350 352 353 354 355 356 357 358 360 361 362 364 365
+ 367 368 369 370 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387
+ 388 389 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408
+ 409 410 411 412 413 414 415 417 418 419 420 421 422 423 424 425 426 427 428 429
+ 430 431 432 433 434 436 437 438 439 441 442 443 444 446 447 448 449 450 451 452
+ 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472
+ 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492
+ 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512
+ 513 514 515 517 518 519 520 522 523 525 526 527 528 529 530 531 532 533 535 536
+ 537 538 539 540 541 542 543 544 546 547 548 549 550 551 552 553 554 555 556 557
+ 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577
+ 578 580 581 582 583 585 586 587 588 589 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 626 627 629 631 632 633 634 636 637 639 644 645 647 649 650 651
+ 653 654 655 658 659 661 662 664 665 666 667 668 670 672 673 674 675 678 680 682
+ 684 687 690 691 692 693 694 695 696 697 698 699 700 701 704 705 707 709 710 712
+ 713 714 715 718 719 720 721 722 723 724 725 726 727 728 729 730 731 732 733 734
+ 735 736 737 738 739 740 741 742 743 744 745 748 749 750 751 752 753 754 755 756
+ 757 758 759 760 761 762 763 764 765 766 767 768 769 770 772 773 775 776 777 778
+ 779 783 784 786 787 788 789 790 791 792 793 794 796 797 798 799 800 801 803 804
+ 805 806 807 808 809 810 811 812 813 816 819 820 821 832 834 835 837 1758 1759
** N=22275 EP=699 IP=10584 FDC=0
X0 1894 3 1895 1 1915 NAND2X1 $T=710820 1682800 0 180 $X=708840 $Y=1677360
X1 1930 3 1916 1 1917 NAND2X1 $T=715440 1672720 0 180 $X=713460 $Y=1667280
X2 2014 3 54 1 44 NAND2X1 $T=744480 1622320 1 180 $X=742500 $Y=1621918
X3 2007 3 2008 1 1970 NAND2X1 $T=743160 1652560 1 0 $X=743158 $Y=1647120
X4 2057 3 2054 1 2008 NAND2X1 $T=751080 1642480 1 180 $X=749100 $Y=1642078
X5 59 3 2059 1 2005 NAND2X1 $T=755040 1692880 0 180 $X=753060 $Y=1687440
X6 2055 3 2114 1 2068 NAND2X1 $T=772860 1702960 0 0 $X=772858 $Y=1702558
X7 2133 3 2113 1 2112 NAND2X1 $T=781440 1682800 1 0 $X=781438 $Y=1677360
X8 66 3 2144 1 2115 NAND2X1 $T=785400 1753360 0 0 $X=785398 $Y=1752958
X9 2181 3 2171 1 2067 NAND2X1 $T=796620 1642480 0 180 $X=794640 $Y=1637040
X10 2226 3 2217 1 2157 NAND2X1 $T=804540 1662640 1 180 $X=802560 $Y=1662238
X11 2261 3 2245 1 2243 NAND2X1 $T=813120 1743280 1 180 $X=811140 $Y=1742878
X12 2292 3 2261 1 2246 NAND2X1 $T=820380 1743280 1 180 $X=818400 $Y=1742878
X13 2247 3 71 1 2274 NAND2X1 $T=821700 1642480 1 180 $X=819720 $Y=1642078
X14 2312 3 2291 1 2292 NAND2X1 $T=838860 1743280 1 0 $X=838858 $Y=1737840
X15 75 3 2302 1 79 NAND2X1 $T=850740 1773520 0 0 $X=850738 $Y=1773118
X16 2347 3 2352 1 2286 NAND2X1 $T=852720 1763440 1 0 $X=852718 $Y=1758000
X17 99 3 2154 1 2551 NAND2X1 $T=888360 1622320 0 180 $X=886380 $Y=1616880
X18 100 3 2476 1 2533 NAND2X1 $T=896280 1622320 1 180 $X=894300 $Y=1621918
X19 2556 3 2537 1 2536 NAND2X1 $T=903540 1662640 1 180 $X=901560 $Y=1662238
X20 2510 3 2537 1 2571 NAND2X1 $T=906840 1652560 0 0 $X=906838 $Y=1652158
X21 2551 3 2476 1 2585 NAND2X1 $T=912120 1622320 0 0 $X=912118 $Y=1621918
X22 2927 3 2914 1 2915 NAND2X1 $T=1016400 1713040 1 180 $X=1014420 $Y=1712638
X23 143 3 142 1 2897 NAND2X1 $T=1017720 1672720 0 180 $X=1015740 $Y=1667280
X24 2926 3 2880 1 2815 NAND2X1 $T=1019040 1642480 0 180 $X=1017060 $Y=1637040
X25 2898 3 145 1 2926 NAND2X1 $T=1019700 1632400 0 0 $X=1019698 $Y=1631998
X26 2959 3 2914 1 2903 NAND2X1 $T=1026960 1702960 1 180 $X=1024980 $Y=1702558
X27 2958 3 2923 1 147 NAND2X1 $T=1029600 1763440 0 0 $X=1029598 $Y=1763038
X28 151 3 2923 1 2968 NAND2X1 $T=1034880 1763440 1 180 $X=1032900 $Y=1763038
X29 153 3 154 1 2983 NAND2X1 $T=1045440 1692880 1 0 $X=1045438 $Y=1687440
X30 155 3 3005 1 148 NAND2X1 $T=1048080 1773520 0 180 $X=1046100 $Y=1768080
X31 152 3 156 1 2958 NAND2X1 $T=1048080 1753360 0 0 $X=1048078 $Y=1752958
X32 161 3 160 1 2927 NAND2X1 $T=1052700 1713040 0 180 $X=1050720 $Y=1707600
X33 176 3 3118 1 174 NAND2X1 $T=1085700 1773520 0 180 $X=1083720 $Y=1768080
X34 3187 3 3135 1 3192 NAND2X1 $T=1102860 1713040 0 180 $X=1100880 $Y=1707600
X35 3185 3 3162 1 3190 NAND2X1 $T=1102860 1753360 0 180 $X=1100880 $Y=1747920
X36 179 3 186 1 3185 NAND2X1 $T=1103520 1733200 1 0 $X=1103518 $Y=1727760
X37 185 3 179 1 3193 NAND2X1 $T=1111440 1753360 0 0 $X=1111438 $Y=1752958
X38 3244 3 3150 1 3225 NAND2X1 $T=1116720 1713040 0 180 $X=1114740 $Y=1707600
X39 184 3 189 1 3213 NAND2X1 $T=1119360 1652560 0 180 $X=1117380 $Y=1647120
X40 186 3 178 1 3244 NAND2X1 $T=1126620 1702960 1 0 $X=1126618 $Y=1697520
X41 30 3 193 1 3288 NAND2X1 $T=1135860 1723120 0 0 $X=1135858 $Y=1722718
X42 344 3 2743 1 3964 NAND2X1 $T=1346400 1713040 1 0 $X=1346398 $Y=1707600
X43 3964 3 4007 1 4030 NAND2X1 $T=1364880 1713040 1 0 $X=1364878 $Y=1707600
X44 4026 3 4029 1 4010 NAND2X1 $T=1368840 1662640 0 0 $X=1368838 $Y=1662238
X45 353 3 2620 1 4060 NAND2X1 $T=1376100 1622320 1 180 $X=1374120 $Y=1621918
X46 4060 3 4077 1 360 NAND2X1 $T=1388640 1622320 1 0 $X=1388638 $Y=1616880
X47 367 3 368 1 369 NAND2X1 $T=1419660 1622320 1 0 $X=1419658 $Y=1616880
X48 4378 3 393 1 4380 NAND2X1 $T=1471140 1753360 0 180 $X=1469160 $Y=1747920
X49 4567 3 413 1 4529 NAND2X1 $T=1521300 1773520 0 180 $X=1519320 $Y=1768080
X50 4633 3 4628 1 4601 NAND2X1 $T=1549680 1692880 0 180 $X=1547700 $Y=1687440
X51 4662 3 413 1 434 NAND2X1 $T=1555620 1773520 0 0 $X=1555618 $Y=1773118
X52 4706 3 4702 1 4628 NAND2X1 $T=1569480 1702960 1 180 $X=1567500 $Y=1702558
X53 437 3 429 1 4714 NAND2X1 $T=1571460 1622320 1 0 $X=1571458 $Y=1616880
X54 4436 3 4748 1 4757 NAND2X1 $T=1580700 1753360 1 0 $X=1580698 $Y=1747920
X55 421 3 4757 1 4753 NAND2X1 $T=1584000 1753360 1 0 $X=1583998 $Y=1747920
X56 455 3 4730 1 4852 NAND2X1 $T=1604460 1672720 1 0 $X=1604458 $Y=1667280
X57 456 3 4849 1 4853 NAND2X1 $T=1606440 1672720 1 0 $X=1606438 $Y=1667280
X58 4936 3 4917 1 5010 NAND2X1 $T=1636140 1702960 1 180 $X=1634160 $Y=1702558
X59 4963 3 4959 1 466 NAND2X1 $T=1645380 1773520 1 180 $X=1643400 $Y=1773118
X60 4946 3 4975 1 4979 NAND2X1 $T=1647360 1702960 1 0 $X=1647358 $Y=1697520
X61 4985 3 4975 1 4963 NAND2X1 $T=1649340 1763440 0 180 $X=1647360 $Y=1758000
X62 5008 3 422 1 5012 NAND2X1 $T=1652640 1723120 1 0 $X=1652638 $Y=1717680
X63 5049 3 422 1 5009 NAND2X1 $T=1665180 1713040 0 180 $X=1663200 $Y=1707600
X64 5259 3 5246 1 5229 NAND2X1 $T=1739760 1692880 1 180 $X=1737780 $Y=1692478
X65 5313 3 5302 1 5235 NAND2X1 $T=1755600 1723120 0 180 $X=1753620 $Y=1717680
X66 5332 3 498 1 5335 NAND2X1 $T=1762860 1773520 1 180 $X=1760880 $Y=1773118
X67 5346 3 5371 1 5359 NAND2X1 $T=1778040 1662640 1 0 $X=1778038 $Y=1657200
X68 5383 3 511 1 5373 NAND2X1 $T=1784640 1743280 0 180 $X=1782660 $Y=1737840
X69 504 3 508 1 5390 NAND2X1 $T=1785960 1702960 0 0 $X=1785958 $Y=1702558
X70 5464 3 5406 1 5418 NAND2X1 $T=1793220 1662640 1 180 $X=1791240 $Y=1662238
X71 362 3 497 1 5456 NAND2X1 $T=1800480 1622320 1 180 $X=1798500 $Y=1621918
X72 5501 3 539 1 5506 NAND2X1 $T=1822260 1773520 1 180 $X=1820280 $Y=1773118
X73 5609 3 5488 1 5478 NAND2X1 $T=1826880 1733200 0 180 $X=1824900 $Y=1727760
X74 5516 3 5509 1 5514 NAND2X1 $T=1828200 1713040 0 180 $X=1826220 $Y=1707600
X75 508 3 586 1 5503 NAND2X1 $T=1841400 1753360 1 0 $X=1841398 $Y=1747920
X76 5541 3 553 1 5550 NAND2X1 $T=1844040 1743280 0 180 $X=1842060 $Y=1737840
X77 576 3 509 1 5595 NAND2X1 $T=1857240 1753360 1 180 $X=1855260 $Y=1752958
X78 5729 3 5551 1 5616 NAND2X1 $T=1887600 1733200 1 180 $X=1885620 $Y=1732798
X79 6032 3 622 1 627 NAND2X1 $T=2003100 1642480 0 0 $X=2003098 $Y=1642078
X80 6257 3 653 1 6212 NAND2X1 $T=2088900 1702960 0 180 $X=2086920 $Y=1697520
X81 6250 3 6268 1 6259 NAND2X1 $T=2089560 1642480 1 0 $X=2089558 $Y=1637040
X82 6246 3 655 1 6213 NAND2X1 $T=2094840 1723120 0 0 $X=2094838 $Y=1722718
X83 6291 3 658 1 6325 NAND2X1 $T=2100120 1632400 1 0 $X=2100118 $Y=1626960
X84 6357 3 6358 1 6354 NAND2X1 $T=2111340 1682800 1 0 $X=2111338 $Y=1677360
X85 6341 3 661 1 6255 NAND2X1 $T=2113980 1642480 0 0 $X=2113978 $Y=1642078
X86 667 3 664 1 6357 NAND2X1 $T=2119920 1672720 0 180 $X=2117940 $Y=1667280
X87 6366 3 6372 1 6404 NAND2X1 $T=2128500 1713040 0 0 $X=2128498 $Y=1712638
X88 6401 3 6459 1 6442 NAND2X1 $T=2144340 1713040 0 0 $X=2144338 $Y=1712638
X89 6505 3 6471 1 6478 NAND2X1 $T=2148960 1672720 0 180 $X=2146980 $Y=1667280
X90 673 3 678 1 6436 NAND2X1 $T=2150940 1632400 1 0 $X=2150938 $Y=1626960
X91 680 3 674 1 6399 NAND2X1 $T=2154240 1622320 0 180 $X=2152260 $Y=1616880
X92 6503 3 6519 1 6505 NAND2X1 $T=2158200 1682800 1 180 $X=2156220 $Y=1682398
X93 6567 3 6546 1 6562 NAND2X1 $T=2177340 1652560 1 180 $X=2175360 $Y=1652158
X94 6547 3 6564 1 6566 NAND2X1 $T=2183280 1682800 0 0 $X=2183278 $Y=1682398
X95 6617 3 6567 1 6552 NAND2X1 $T=2190540 1652560 1 180 $X=2188560 $Y=1652158
X96 6710 3 6728 1 6724 NAND2X1 $T=2220240 1652560 0 0 $X=2220238 $Y=1652158
X97 6712 3 6747 1 6748 NAND2X1 $T=2225520 1713040 1 0 $X=2225518 $Y=1707600
X98 6747 3 6799 1 6782 NAND2X1 $T=2248620 1713040 1 0 $X=2248618 $Y=1707600
X99 6855 3 704 1 6843 NAND2X1 $T=2263140 1773520 1 0 $X=2263138 $Y=1768080
X100 6874 3 6891 1 6781 NAND2X1 $T=2269080 1652560 1 0 $X=2269078 $Y=1647120
X101 6907 3 6909 1 6937 NAND2X1 $T=2277660 1713040 1 0 $X=2277658 $Y=1707600
X102 6932 3 6959 1 6945 NAND2X1 $T=2291520 1692880 0 0 $X=2291518 $Y=1692478
X103 6928 3 6938 1 719 NAND2X1 $T=2304060 1632400 1 0 $X=2304058 $Y=1626960
X104 7029 3 7040 1 721 NAND2X1 $T=2310660 1632400 1 0 $X=2310658 $Y=1626960
X105 7045 3 7086 1 7065 NAND2X1 $T=2329800 1682800 0 0 $X=2329798 $Y=1682398
X106 7070 3 726 1 733 NAND2X1 $T=2335080 1763440 0 0 $X=2335078 $Y=1763038
X107 772 3 632 1 7633 NAND2X1 $T=2502060 1692880 1 180 $X=2500080 $Y=1692478
X108 772 3 626 1 7777 NAND2X1 $T=2541000 1632400 0 180 $X=2539020 $Y=1626960
X109 8045 3 805 1 808 NAND2X1 $T=2608980 1632400 0 180 $X=2607000 $Y=1626960
X110 7925 3 7948 1 8074 NAND2X1 $T=2609640 1662640 1 0 $X=2609638 $Y=1657200
X111 8095 3 7963 1 8054 NAND2X1 $T=2618220 1702960 0 180 $X=2616240 $Y=1697520
X112 8056 3 8073 1 8047 NAND2X1 $T=2621520 1672720 1 0 $X=2621518 $Y=1667280
X113 1894 1 3 1895 1896 NOR2X4 $T=710160 1672720 0 180 $X=705540 $Y=1667280
X114 59 1 3 2059 2080 NOR2X4 $T=757020 1692880 1 0 $X=757018 $Y=1687440
X115 3770 1 3 3842 3844 NOR2X4 $T=1302840 1632400 1 180 $X=1298220 $Y=1631998
X116 3842 1 3 316 283 NOR2X4 $T=1304820 1652560 1 0 $X=1304818 $Y=1647120
X117 3842 1 3 316 226 NOR2X4 $T=1309440 1662640 1 180 $X=1304820 $Y=1662238
X118 316 1 3 4460 4463 NOR2X4 $T=1497540 1632400 1 180 $X=1492920 $Y=1631998
X119 399 1 3 400 4501 NOR2X4 $T=1501500 1642480 0 0 $X=1501498 $Y=1642078
X120 395 1 3 4501 407 NOR2X4 $T=1506120 1642480 0 0 $X=1506118 $Y=1642078
X121 4514 1 3 4512 4524 NOR2X4 $T=1514040 1713040 0 180 $X=1509420 $Y=1707600
X122 415 1 3 4552 4572 NOR2X4 $T=1522620 1702960 1 0 $X=1522618 $Y=1697520
X123 316 1 3 424 4581 NOR2X4 $T=1544400 1662640 0 180 $X=1539780 $Y=1657200
X124 406 1 3 424 429 NOR2X4 $T=1554960 1632400 0 180 $X=1550340 $Y=1626960
X125 431 1 3 4685 415 NOR2X4 $T=1558920 1692880 1 0 $X=1558918 $Y=1687440
X126 427 1 3 4721 4706 NOR2X4 $T=1578720 1702960 1 180 $X=1574100 $Y=1702558
X127 427 1 3 4721 4755 NOR2X4 $T=1586640 1702960 1 180 $X=1582020 $Y=1702558
X128 406 1 3 424 4765 NOR2X4 $T=1589940 1662640 1 0 $X=1589938 $Y=1657200
X129 4785 1 3 4779 4799 NOR2X4 $T=1593240 1713040 0 0 $X=1593238 $Y=1712638
X130 4798 1 3 4779 4742 NOR2X4 $T=1595220 1702960 1 0 $X=1595218 $Y=1697520
X131 4832 1 3 4755 4857 NOR2X4 $T=1609740 1743280 1 0 $X=1609738 $Y=1737840
X132 4849 1 3 4895 4887 NOR2X4 $T=1620960 1743280 1 0 $X=1620958 $Y=1737840
X133 316 1 3 5303 493 NOR2X4 $T=1769460 1632400 1 180 $X=1764840 $Y=1631998
X134 6032 1 3 622 624 NOR2X4 $T=1999800 1642480 1 180 $X=1995180 $Y=1642078
X135 47 3 44 1927 1 NAND2BX1 $T=718740 1622320 1 180 $X=716100 $Y=1621918
X136 42 3 41 1953 1 NAND2BX1 $T=717420 1773520 1 0 $X=717418 $Y=1768080
X137 2103 3 2067 2057 1 NAND2BX1 $T=757680 1642480 1 180 $X=755040 $Y=1642078
X138 2116 3 2115 2168 1 NAND2BX1 $T=786720 1743280 0 0 $X=786718 $Y=1742878
X139 2152 3 2157 2084 1 NAND2BX1 $T=792000 1672720 0 180 $X=789360 $Y=1667280
X140 2279 3 2286 72 1 NAND2BX1 $T=826980 1763440 1 180 $X=824340 $Y=1763038
X141 2912 3 2897 2862 1 NAND2BX1 $T=1012440 1682800 1 180 $X=1009800 $Y=1682398
X142 3186 3 3152 3164 1 NAND2BX1 $T=1100220 1642480 1 180 $X=1097580 $Y=1642078
X143 3216 3 3213 3211 1 NAND2BX1 $T=1118700 1662640 0 0 $X=1118698 $Y=1662238
X144 4572 3 380 4599 1 NAND2BX1 $T=1531860 1692880 1 0 $X=1531858 $Y=1687440
X145 4747 3 421 4752 1 NAND2BX1 $T=1581360 1743280 1 0 $X=1581358 $Y=1737840
X146 451 3 4625 4748 1 NAND2BX1 $T=1584000 1773520 0 180 $X=1581360 $Y=1768080
X147 4514 3 4773 4781 1 NAND2BX1 $T=1590600 1743280 0 0 $X=1590598 $Y=1742878
X148 4702 3 4911 4929 1 NAND2BX1 $T=1624920 1753360 0 0 $X=1624918 $Y=1752958
X149 487 3 5301 5311 1 NAND2BX1 $T=1751640 1672720 0 0 $X=1751638 $Y=1672318
X150 6110 3 6112 6098 1 NAND2BX1 $T=2052600 1753360 1 180 $X=2049960 $Y=1752958
X151 6223 3 6213 6182 1 NAND2BX1 $T=2077020 1733200 1 180 $X=2074380 $Y=1732798
X152 6563 3 6566 6479 1 NAND2BX1 $T=2178000 1662640 0 180 $X=2175360 $Y=1657200
X153 6728 3 6731 6727 1 NAND2BX1 $T=2222220 1642480 0 0 $X=2222218 $Y=1642078
X154 6772 3 6729 6754 1 NAND2BX1 $T=2230140 1672720 0 180 $X=2227500 $Y=1667280
X155 6858 3 6843 6901 1 NAND2BX1 $T=2269740 1743280 1 0 $X=2269738 $Y=1737840
X156 7634 3 7633 7637 1 NAND2BX1 $T=2507340 1713040 1 0 $X=2507338 $Y=1707600
X157 1930 1896 3 1915 1 1929 OAI21X1 $T=719400 1682800 0 180 $X=716100 $Y=1677360
X158 2103 2117 3 2067 1 2121 OAI21X1 $T=775500 1642480 1 0 $X=775498 $Y=1637040
X159 2912 2913 3 2897 1 2869 OAI21X1 $T=1015740 1692880 1 180 $X=1012440 $Y=1692478
X160 2945 2900 3 2927 1 2946 OAI21X1 $T=1025640 1713040 0 0 $X=1025638 $Y=1712638
X161 2968 149 3 2919 1 2966 OAI21X1 $T=1034220 1753360 1 180 $X=1030920 $Y=1752958
X162 4275 383 3 384 1 4264 OAI21X1 $T=1449360 1773520 0 0 $X=1449358 $Y=1773118
X163 4977 4986 3 5012 1 5005 OAI21X1 $T=1654620 1723120 1 0 $X=1654618 $Y=1717680
X164 6183 6223 3 6213 1 6215 OAI21X1 $T=2076360 1733200 0 180 $X=2073060 $Y=1727760
X165 6562 6521 3 6576 1 692 OAI21X1 $T=2175360 1652560 1 0 $X=2175358 $Y=1647120
X166 5921 5920 3 7119 1 7123 OAI21X1 $T=2344980 1733200 0 0 $X=2344978 $Y=1732798
X167 2118 3 2094 2112 1 2083 OAI21XL $T=770220 1672720 0 180 $X=767580 $Y=1667280
X168 2105 3 2094 2117 1 2054 OAI21XL $T=774840 1652560 0 180 $X=772200 $Y=1647120
X169 2112 3 2152 2157 1 2216 OAI21XL $T=799260 1672720 1 0 $X=799258 $Y=1667280
X170 79 3 2279 2286 1 2258 OAI21XL $T=832920 1763440 0 0 $X=832918 $Y=1763038
X171 2382 3 104 2550 1 2588 OAI21XL $T=906840 1713040 1 0 $X=906838 $Y=1707600
X172 2903 3 2900 2913 1 2830 OAI21XL $T=1015080 1713040 0 180 $X=1012440 $Y=1707600
X173 3216 3 3197 3213 1 3120 OAI21XL $T=1106820 1662640 1 180 $X=1104180 $Y=1662238
X174 3963 3 3894 3954 1 3936 OAI21XL $T=1342440 1682800 0 180 $X=1339800 $Y=1677360
X175 399 3 4472 397 1 4335 OAI21XL $T=1494240 1662640 1 180 $X=1491600 $Y=1662238
X176 4752 3 4706 4753 1 4749 OAI21XL $T=1582680 1733200 1 0 $X=1582678 $Y=1727760
X177 444 3 455 446 1 4837 OAI21XL $T=1607760 1622320 1 0 $X=1607758 $Y=1616880
X178 6110 3 639 6112 1 6115 OAI21XL $T=2042040 1753360 0 0 $X=2042038 $Y=1752958
X179 6400 3 6403 6404 1 6409 OAI21XL $T=2127180 1702960 1 0 $X=2127178 $Y=1697520
X180 6404 3 6435 6442 1 6441 OAI21XL $T=2139060 1713040 1 0 $X=2139058 $Y=1707600
X181 5814 3 602 6523 1 682 OAI21XL $T=2159520 1753360 0 0 $X=2159518 $Y=1752958
X182 668 3 6342 623 1 6523 OAI21XL $T=2167440 1753360 1 180 $X=2164800 $Y=1752958
X183 6505 3 6563 6566 1 6549 OAI21XL $T=2176680 1672720 1 0 $X=2176678 $Y=1667280
X184 6622 3 6637 6680 1 690 OAI21XL $T=2205720 1773520 1 0 $X=2205718 $Y=1768080
X185 6712 3 6684 6705 1 6711 OAI21XL $T=2219580 1702960 1 180 $X=2216940 $Y=1702558
X186 6772 3 6764 6729 1 6784 OAI21XL $T=2234100 1672720 0 0 $X=2234098 $Y=1672318
X187 6785 3 695 6764 1 6766 OAI21XL $T=2236740 1692880 0 180 $X=2234100 $Y=1687440
X188 6782 3 695 6773 1 6706 OAI21XL $T=2236740 1713040 0 180 $X=2234100 $Y=1707600
X189 6786 3 698 6781 1 6780 OAI21XL $T=2238060 1632400 0 180 $X=2235420 $Y=1626960
X190 6844 3 6843 6842 1 6767 OAI21XL $T=2252580 1743280 0 180 $X=2249940 $Y=1737840
X191 6857 3 695 6856 1 6859 OAI21XL $T=2256540 1672720 0 0 $X=2256538 $Y=1672318
X192 6872 3 695 6870 1 6871 OAI21XL $T=2263140 1723120 0 180 $X=2260500 $Y=1717680
X193 6857 3 695 6889 1 707 OAI21XL $T=2268420 1672720 0 0 $X=2268418 $Y=1672318
X194 6858 3 695 6843 1 6908 OAI21XL $T=2269740 1753360 1 0 $X=2269738 $Y=1747920
X195 623 3 621 6353 1 6977 OAI21XL $T=2288880 1733200 1 0 $X=2288878 $Y=1727760
X196 714 3 7014 6937 1 7022 OAI21XL $T=2299440 1713040 1 0 $X=2299438 $Y=1707600
X197 7023 3 5814 7049 1 7050 OAI21XL $T=2315280 1753360 1 0 $X=2315278 $Y=1747920
X198 7123 3 602 7160 1 7151 OAI21XL $T=2356860 1733200 0 0 $X=2356858 $Y=1732798
X199 633 3 623 727 1 7119 OAI21XL $T=2384580 1733200 0 0 $X=2384578 $Y=1732798
X200 7222 3 7248 7250 1 7249 OAI21XL $T=2388540 1692880 0 0 $X=2388538 $Y=1692478
X201 7301 3 7260 727 1 7257 OAI21XL $T=2396460 1753360 0 180 $X=2393820 $Y=1747920
X202 5921 3 718 7313 1 7314 OAI21XL $T=2407020 1702960 1 0 $X=2407018 $Y=1697520
X203 623 3 605 7314 1 751 OAI21XL $T=2407020 1702960 0 0 $X=2407018 $Y=1702558
X204 748 3 752 749 1 753 OAI21XL $T=2414940 1773520 0 180 $X=2412300 $Y=1768080
X205 756 3 633 754 1 7348 OAI21XL $T=2420220 1632400 1 180 $X=2417580 $Y=1631998
X206 7331 3 7329 7347 1 7315 OAI21XL $T=2420880 1753360 1 0 $X=2420878 $Y=1747920
X207 5929 3 621 7371 1 7347 OAI21XL $T=2427480 1723120 1 180 $X=2424840 $Y=1722718
X208 668 3 7395 5936 1 7403 OAI21XL $T=2434080 1723120 1 0 $X=2434078 $Y=1717680
X209 607 3 602 7403 1 7411 OAI21XL $T=2435400 1713040 1 0 $X=2435398 $Y=1707600
X210 632 3 631 668 1 7397 OAI21XL $T=2438040 1642480 1 180 $X=2435400 $Y=1642078
X211 614 3 758 727 1 7371 OAI21XL $T=2443320 1723120 1 180 $X=2440680 $Y=1722718
X212 7262 3 610 7397 1 7492 OAI21XL $T=2443320 1652560 1 0 $X=2443318 $Y=1647120
X213 623 3 634 5919 1 7420 OAI21XL $T=2443320 1682800 1 0 $X=2443318 $Y=1677360
X214 7416 3 5921 7420 1 7444 OAI21XL $T=2443320 1692880 1 0 $X=2443318 $Y=1687440
X215 621 3 626 6166 1 7466 OAI21XL $T=2451240 1672720 1 0 $X=2451238 $Y=1667280
X216 7313 3 758 632 1 7493 OAI21XL $T=2459160 1723120 0 0 $X=2459158 $Y=1722718
X217 7492 3 7491 7494 1 7510 OAI21XL $T=2463120 1682800 1 0 $X=2463118 $Y=1677360
X218 631 3 758 6342 1 7527 OAI21XL $T=2465760 1702960 0 0 $X=2465758 $Y=1702558
X219 7479 3 7511 7537 1 765 OAI21XL $T=2481600 1713040 0 0 $X=2481598 $Y=1712638
X220 766 3 758 7580 1 7582 OAI21XL $T=2491500 1652560 0 0 $X=2491498 $Y=1652158
X221 5929 3 768 633 1 7580 OAI21XL $T=2496780 1652560 0 0 $X=2496778 $Y=1652158
X222 7587 3 7556 7444 1 7638 OAI21XL $T=2496780 1743280 1 0 $X=2496778 $Y=1737840
X223 7634 3 614 7633 1 7587 OAI21XL $T=2502060 1713040 0 180 $X=2499420 $Y=1707600
X224 7635 3 7636 7641 1 7644 OAI21XL $T=2503380 1642480 1 0 $X=2503378 $Y=1637040
X225 7262 3 776 756 1 7675 OAI21XL $T=2508660 1662640 0 0 $X=2508658 $Y=1662238
X226 7634 3 776 7633 1 7703 OAI21XL $T=2508660 1692880 1 0 $X=2508658 $Y=1687440
X227 776 3 768 727 1 7676 OAI21XL $T=2513940 1723120 0 180 $X=2511300 $Y=1717680
X228 626 3 772 623 1 7718 OAI21XL $T=2515260 1642480 0 0 $X=2515258 $Y=1642078
X229 778 3 631 7675 1 7697 OAI21XL $T=2515260 1662640 0 0 $X=2515258 $Y=1662238
X230 607 3 763 754 1 7684 OAI21XL $T=2517900 1622320 0 180 $X=2515260 $Y=1616880
X231 7721 3 7719 7730 1 7815 OAI21XL $T=2536380 1763440 0 0 $X=2536378 $Y=1763038
X232 634 3 626 633 1 7803 OAI21XL $T=2537700 1642480 0 0 $X=2537698 $Y=1642078
X233 600 3 772 7684 1 7783 OAI21XL $T=2541660 1622320 0 180 $X=2539020 $Y=1616880
X234 786 3 7550 631 1 7825 OAI21XL $T=2544960 1702960 0 0 $X=2544958 $Y=1702558
X235 7818 3 7733 7827 1 7862 OAI21XL $T=2546940 1723120 0 0 $X=2546938 $Y=1722718
X236 7804 3 7800 7837 1 7827 OAI21XL $T=2549580 1682800 1 0 $X=2549578 $Y=1677360
X237 7836 3 7801 7815 1 7816 OAI21XL $T=2552220 1763440 1 180 $X=2549580 $Y=1763038
X238 7703 3 7701 794 1 7900 OAI21XL $T=2568720 1652560 0 0 $X=2568718 $Y=1652158
X239 7825 3 7781 7887 1 7928 OAI21XL $T=2568720 1692880 1 0 $X=2568718 $Y=1687440
X240 7912 3 7465 7783 1 7916 OAI21XL $T=2577960 1733200 0 0 $X=2577958 $Y=1732798
X241 797 3 7931 7941 1 7944 OAI21XL $T=2584560 1753360 1 180 $X=2581920 $Y=1752958
X242 803 3 7509 7495 1 7990 OAI21XL $T=2600400 1733200 1 180 $X=2597760 $Y=1732798
X243 8059 3 8086 820 1 8093 OAI21XL $T=2622840 1713040 1 180 $X=2620200 $Y=1712638
X244 2164 2142 2227 3 1 XOR2X4 $T=790680 1702960 0 0 $X=790678 $Y=1702558
X245 6739 6709 691 3 1 XOR2X4 $T=2224860 1622320 0 180 $X=2213640 $Y=1616880
X246 7044 7027 5958 3 1 XOR2X4 $T=2315280 1702960 0 180 $X=2304060 $Y=1697520
X247 1930 3 1 1965 INVX1 $T=719400 1672720 1 0 $X=719398 $Y=1667280
X248 47 3 1 1945 INVX1 $T=726000 1622320 0 180 $X=724680 $Y=1616880
X249 1963 3 1 1964 INVX1 $T=730620 1713040 1 180 $X=729300 $Y=1712638
X250 1981 3 1 1916 INVX1 $T=737220 1682800 1 0 $X=737218 $Y=1677360
X251 63 3 1 65 INVX1 $T=766260 1773520 0 0 $X=766258 $Y=1773118
X252 2068 3 1 2140 INVX1 $T=777480 1702960 0 0 $X=777478 $Y=1702558
X253 2085 3 1 2137 INVX1 $T=780120 1713040 0 0 $X=780118 $Y=1712638
X254 64 3 1 2150 INVX1 $T=782100 1773520 0 0 $X=782098 $Y=1773118
X255 2216 3 1 2117 INVX1 $T=784080 1662640 0 180 $X=782760 $Y=1657200
X256 69 3 1 70 INVX1 $T=811800 1773520 0 180 $X=810480 $Y=1768080
X257 2292 3 1 2262 INVX1 $T=830280 1743280 0 180 $X=828960 $Y=1737840
X258 2494 3 1 2537 INVX1 $T=898920 1662640 0 0 $X=898918 $Y=1662238
X259 37 3 1 2509 INVX1 $T=903540 1753360 0 180 $X=902220 $Y=1747920
X260 2551 3 1 105 INVX1 $T=907500 1622320 1 0 $X=907498 $Y=1616880
X261 2516 3 1 2556 INVX1 $T=911460 1672720 1 180 $X=910140 $Y=1672318
X262 2588 3 1 2579 INVX1 $T=920700 1723120 0 0 $X=920698 $Y=1722718
X263 28 3 1 2576 INVX1 $T=933900 1652560 1 0 $X=933898 $Y=1647120
X264 103 3 1 2614 INVX1 $T=933900 1682800 0 0 $X=933898 $Y=1682398
X265 30 3 1 2542 INVX1 $T=974160 1733200 0 180 $X=972840 $Y=1727760
X266 137 3 1 2805 INVX1 $T=999240 1642480 0 0 $X=999238 $Y=1642078
X267 2945 3 1 2914 INVX1 $T=1021020 1713040 1 180 $X=1019700 $Y=1712638
X268 2926 3 1 2883 INVX1 $T=1021680 1642480 0 180 $X=1020360 $Y=1637040
X269 2958 3 1 2922 INVX1 $T=1023660 1763440 0 180 $X=1022340 $Y=1758000
X270 148 3 1 2925 INVX1 $T=1024980 1773520 1 180 $X=1023660 $Y=1773118
X271 2983 3 1 2988 INVX1 $T=1039500 1702960 0 180 $X=1038180 $Y=1697520
X272 2927 3 1 2986 INVX1 $T=1047420 1713040 0 180 $X=1046100 $Y=1707600
X273 163 3 1 164 INVX1 $T=1059300 1743280 0 0 $X=1059298 $Y=1742878
X274 174 3 1 170 INVX1 $T=1077120 1773520 1 180 $X=1075800 $Y=1773118
X275 3167 3 1 3197 INVX1 $T=1098240 1672720 1 0 $X=1098238 $Y=1667280
X276 3193 3 1 3172 INVX1 $T=1102200 1753360 1 180 $X=1100880 $Y=1752958
X277 3187 3 1 3203 INVX1 $T=1103520 1702960 1 0 $X=1103518 $Y=1697520
X278 3244 3 1 3214 INVX1 $T=1120680 1702960 1 180 $X=1119360 $Y=1702558
X279 29 3 1 3297 INVX1 $T=1129920 1632400 1 0 $X=1129918 $Y=1626960
X280 104 3 1 3448 INVX1 $T=1171500 1702960 0 0 $X=1171498 $Y=1702558
X281 184 3 1 3743 INVX1 $T=1270500 1702960 1 0 $X=1270498 $Y=1697520
X282 3964 3 1 4020 INVX1 $T=1354980 1702960 0 0 $X=1354978 $Y=1702558
X283 349 3 1 4025 INVX1 $T=1360260 1642480 0 0 $X=1360258 $Y=1642078
X284 4060 3 1 4096 INVX1 $T=1388640 1632400 1 0 $X=1388638 $Y=1626960
X285 4117 3 1 4092 INVX1 $T=1396560 1642480 1 0 $X=1396558 $Y=1637040
X286 4088 3 1 4131 INVX1 $T=1396560 1652560 1 0 $X=1396558 $Y=1647120
X287 3770 3 1 362 INVX1 $T=1403820 1672720 1 0 $X=1403818 $Y=1667280
X288 373 3 1 4241 INVX1 $T=1428240 1662640 1 0 $X=1428238 $Y=1657200
X289 381 3 1 3868 INVX1 $T=1444740 1642480 0 180 $X=1443420 $Y=1637040
X290 4400 3 1 4272 INVX1 $T=1455300 1733200 1 180 $X=1453980 $Y=1732798
X291 387 3 1 395 INVX1 $T=1461240 1662640 0 0 $X=1461238 $Y=1662238
X292 122 3 1 4365 INVX1 $T=1467180 1733200 1 0 $X=1467178 $Y=1727760
X293 157 3 1 4415 INVX1 $T=1477740 1723120 0 0 $X=1477738 $Y=1722718
X294 4403 3 1 4396 INVX1 $T=1486320 1733200 0 180 $X=1485000 $Y=1727760
X295 4424 3 1 4418 INVX1 $T=1490940 1773520 1 180 $X=1489620 $Y=1773118
X296 130 3 1 405 INVX1 $T=1500180 1773520 1 180 $X=1498860 $Y=1773118
X297 4529 3 1 414 INVX1 $T=1521960 1773520 0 0 $X=1521958 $Y=1773118
X298 4567 3 1 4570 INVX1 $T=1527240 1733200 0 0 $X=1527238 $Y=1732798
X299 380 3 1 4633 INVX1 $T=1548360 1682800 0 0 $X=1548358 $Y=1682398
X300 4714 3 1 4400 INVX1 $T=1559580 1662640 0 180 $X=1558260 $Y=1657200
X301 4586 3 1 4662 INVX1 $T=1560240 1763440 0 180 $X=1558920 $Y=1758000
X302 4528 3 1 425 INVX1 $T=1564200 1733200 1 0 $X=1564198 $Y=1727760
X303 4625 3 1 4692 INVX1 $T=1568160 1763440 1 180 $X=1566840 $Y=1763038
X304 438 3 1 4660 INVX1 $T=1573440 1652560 1 180 $X=1572120 $Y=1652158
X305 4729 3 1 4725 INVX1 $T=1576740 1642480 0 180 $X=1575420 $Y=1637040
X306 4730 3 1 4738 INVX1 $T=1576740 1642480 0 0 $X=1576738 $Y=1642078
X307 428 3 1 4767 INVX1 $T=1591920 1763440 0 0 $X=1591918 $Y=1763038
X308 406 3 1 426 INVX1 $T=1597860 1652560 0 0 $X=1597858 $Y=1652158
X309 4514 3 1 4836 INVX1 $T=1605780 1743280 1 180 $X=1604460 $Y=1742878
X310 4851 3 1 4871 INVX1 $T=1608420 1753360 0 0 $X=1608418 $Y=1752958
X311 4799 3 1 4890 INVX1 $T=1618320 1733200 1 0 $X=1618318 $Y=1727760
X312 4886 3 1 4904 INVX1 $T=1625580 1713040 0 180 $X=1624260 $Y=1707600
X313 4857 3 1 4959 INVX1 $T=1629540 1773520 0 0 $X=1629538 $Y=1773118
X314 463 3 1 3770 INVX1 $T=1636140 1622320 1 180 $X=1634820 $Y=1621918
X315 4946 3 1 4936 INVX1 $T=1636140 1702960 0 180 $X=1634820 $Y=1697520
X316 464 3 1 4971 INVX1 $T=1644720 1763440 0 0 $X=1644718 $Y=1763038
X317 4799 3 1 4975 INVX1 $T=1647360 1723120 0 0 $X=1647358 $Y=1722718
X318 4949 3 1 4977 INVX1 $T=1648020 1723120 1 0 $X=1648018 $Y=1717680
X319 4917 3 1 4986 INVX1 $T=1649340 1723120 1 0 $X=1649338 $Y=1717680
X320 472 3 1 5053 INVX1 $T=1661880 1662640 0 0 $X=1661878 $Y=1662238
X321 457 3 1 4911 INVX1 $T=1672440 1753360 0 0 $X=1672438 $Y=1752958
X322 465 3 1 5070 INVX1 $T=1696200 1692880 1 180 $X=1694880 $Y=1692478
X323 169 3 1 5202 INVX1 $T=1720620 1763440 0 0 $X=1720618 $Y=1763038
X324 5202 3 1 5203 INVX1 $T=1723260 1763440 1 0 $X=1723258 $Y=1758000
X325 251 3 1 5301 INVX1 $T=1740420 1672720 1 0 $X=1740418 $Y=1667280
X326 272 3 1 5280 INVX1 $T=1752960 1743280 1 0 $X=1752958 $Y=1737840
X327 507 3 1 496 INVX1 $T=1777380 1733200 0 180 $X=1776060 $Y=1727760
X328 517 3 1 504 INVX1 $T=1789920 1682800 0 180 $X=1788600 $Y=1677360
X329 543 3 1 546 INVX1 $T=1833480 1622320 0 0 $X=1833478 $Y=1621918
X330 5548 3 1 5534 INVX1 $T=1840080 1773520 0 180 $X=1838760 $Y=1768080
X331 5757 3 1 5787 INVX1 $T=1928520 1662640 1 0 $X=1928518 $Y=1657200
X332 6115 3 1 6183 INVX1 $T=2044680 1743280 0 0 $X=2044678 $Y=1742878
X333 6214 3 1 6181 INVX1 $T=2071080 1753360 1 180 $X=2069760 $Y=1752958
X334 6212 3 1 6219 INVX1 $T=2073720 1702960 1 0 $X=2073718 $Y=1697520
X335 6218 3 1 6256 INVX1 $T=2076360 1662640 1 0 $X=2076358 $Y=1657200
X336 6245 3 1 6223 INVX1 $T=2084280 1733200 1 0 $X=2084278 $Y=1727760
X337 6255 3 1 6261 INVX1 $T=2091540 1642480 1 180 $X=2090220 $Y=1642078
X338 6360 3 1 6246 INVX1 $T=2096160 1723120 0 180 $X=2094840 $Y=1717680
X339 6325 3 1 6269 INVX1 $T=2098800 1632400 1 180 $X=2097480 $Y=1631998
X340 6323 3 1 6257 INVX1 $T=2100120 1702960 0 180 $X=2098800 $Y=1697520
X341 6357 3 1 6364 INVX1 $T=2110680 1672720 1 0 $X=2110678 $Y=1667280
X342 6326 3 1 6403 INVX1 $T=2126520 1692880 1 0 $X=2126518 $Y=1687440
X343 6410 3 1 6291 INVX1 $T=2130480 1652560 1 180 $X=2129160 $Y=1652158
X344 6436 3 1 6389 INVX1 $T=2138400 1622320 1 180 $X=2137080 $Y=1621918
X345 6452 3 1 6341 INVX1 $T=2143020 1642480 1 180 $X=2141700 $Y=1642078
X346 6521 3 1 6470 INVX1 $T=2160180 1652560 1 0 $X=2160178 $Y=1647120
X347 6544 3 1 684 INVX1 $T=2168760 1622320 0 180 $X=2167440 $Y=1616880
X348 6617 3 1 6593 INVX1 $T=2195820 1652560 1 180 $X=2194500 $Y=1652158
X349 6710 3 1 6731 INVX1 $T=2217600 1642480 0 0 $X=2217598 $Y=1642078
X350 6781 3 1 6734 INVX1 $T=2237400 1642480 0 180 $X=2236080 $Y=1637040
X351 6775 3 1 6786 INVX1 $T=2245320 1632400 0 180 $X=2244000 $Y=1626960
X352 6784 3 1 6856 INVX1 $T=2257200 1672720 1 0 $X=2257198 $Y=1667280
X353 6799 3 1 6872 INVX1 $T=2261160 1723120 0 0 $X=2261158 $Y=1722718
X354 631 3 1 5900 INVX1 $T=2275020 1652560 0 0 $X=2275018 $Y=1652158
X355 712 3 1 6980 INVX1 $T=2290860 1763440 1 0 $X=2290858 $Y=1758000
X356 6932 3 1 7014 INVX1 $T=2293500 1713040 1 0 $X=2293498 $Y=1707600
X357 714 3 1 7015 INVX1 $T=2311980 1763440 0 0 $X=2311978 $Y=1763038
X358 5936 3 1 7026 INVX1 $T=2318580 1662640 1 180 $X=2317260 $Y=1662238
X359 6959 3 1 7043 INVX1 $T=2319240 1692880 0 0 $X=2319238 $Y=1692478
X360 7065 3 1 7017 INVX1 $T=2321220 1692880 0 180 $X=2319900 $Y=1687440
X361 5919 3 1 7088 INVX1 $T=2350260 1632400 0 180 $X=2348940 $Y=1626960
X362 5929 3 1 7171 INVX1 $T=2356200 1662640 0 0 $X=2356198 $Y=1662238
X363 5936 3 1 7187 INVX1 $T=2366760 1692880 0 0 $X=2366758 $Y=1692478
X364 7327 3 1 740 INVX1 $T=2387220 1773520 1 180 $X=2385900 $Y=1773118
X365 742 3 1 752 INVX1 $T=2401080 1773520 1 0 $X=2401078 $Y=1768080
X366 5919 3 1 7313 INVX1 $T=2408340 1682800 1 0 $X=2408338 $Y=1677360
X367 607 3 1 7395 INVX1 $T=2442660 1713040 1 0 $X=2442658 $Y=1707600
X368 634 3 1 7416 INVX1 $T=2450580 1682800 1 0 $X=2450578 $Y=1677360
X369 7981 3 1 7975 INVX1 $T=2599080 1682800 0 180 $X=2597760 $Y=1677360
X370 799 3 1 8024 INVX1 $T=2600400 1773520 0 0 $X=2600398 $Y=1773118
X371 7980 3 1 8075 INVX1 $T=2613600 1672720 0 0 $X=2613598 $Y=1672318
X372 8054 3 1 8077 INVX1 $T=2615580 1682800 1 0 $X=2615578 $Y=1677360
X373 8081 3 1 8094 INVX1 $T=2620860 1652560 0 0 $X=2620858 $Y=1652158
X374 8061 3 1 8058 INVX1 $T=2622840 1622320 0 180 $X=2621520 $Y=1616880
X375 1961 1916 1 1965 1969 3 AOI21X2 $T=731940 1672720 1 0 $X=731938 $Y=1667280
X376 2142 2137 1 2140 2139 3 AOI21X2 $T=788700 1713040 1 180 $X=784080 $Y=1712638
X377 2868 2865 1 2869 2781 3 AOI21X2 $T=1001220 1692880 1 0 $X=1001218 $Y=1687440
X378 2986 2959 1 2988 2913 3 AOI21X2 $T=1035540 1702960 0 0 $X=1035538 $Y=1702558
X379 3167 3188 1 3164 182 3 AOI21X2 $T=1104840 1652560 0 180 $X=1100220 $Y=1647120
X380 4570 410 1 4514 4597 3 AOI21X2 $T=1570140 1713040 1 0 $X=1570138 $Y=1707600
X381 674 6389 1 675 672 3 AOI21X2 $T=2141700 1622320 1 0 $X=2141698 $Y=1616880
X382 696 6783 1 6780 6709 3 AOI21X2 $T=2236080 1622320 0 0 $X=2236078 $Y=1621918
X383 696 700 1 701 6841 3 AOI21X2 $T=2251920 1652560 1 180 $X=2247300 $Y=1652158
X384 7028 696 1 7022 7027 3 AOI21X2 $T=2313960 1713040 1 0 $X=2313958 $Y=1707600
X385 1 48 1978 1960 3 NOR2X1 $T=731940 1753360 0 0 $X=731938 $Y=1752958
X386 1 2014 54 47 3 NOR2X1 $T=745800 1622320 0 180 $X=743820 $Y=1616880
X387 1 2103 2105 2107 3 NOR2X1 $T=770880 1642480 1 0 $X=770878 $Y=1637040
X388 1 2133 2113 2118 3 NOR2X1 $T=774840 1682800 1 180 $X=772860 $Y=1682398
X389 1 2055 2114 2085 3 NOR2X1 $T=775500 1713040 0 0 $X=775498 $Y=1712638
X390 1 2181 2171 2103 3 NOR2X1 $T=797940 1642480 1 180 $X=795960 $Y=1642078
X391 1 2226 2217 2152 3 NOR2X1 $T=805200 1672720 0 180 $X=803220 $Y=1667280
X392 1 73 2279 2245 3 NOR2X1 $T=826320 1763440 0 180 $X=824340 $Y=1758000
X393 1 75 2302 73 3 NOR2X1 $T=842820 1773520 1 180 $X=840840 $Y=1773118
X394 1 2347 2352 2279 3 NOR2X1 $T=848760 1763440 1 0 $X=848758 $Y=1758000
X395 1 143 142 2912 3 NOR2X1 $T=1017720 1682800 0 180 $X=1015740 $Y=1677360
X396 1 2912 2903 2868 3 NOR2X1 $T=1019700 1692880 1 0 $X=1019698 $Y=1687440
X397 1 161 160 2945 3 NOR2X1 $T=1055340 1713040 1 180 $X=1053360 $Y=1712638
X398 1 185 183 3210 3 NOR2X1 $T=1102860 1632400 1 0 $X=1102858 $Y=1626960
X399 1 3213 3210 3186 3 NOR2X1 $T=1108140 1642480 0 180 $X=1106160 $Y=1637040
X400 1 3216 3210 3188 3 NOR2X1 $T=1109460 1652560 0 180 $X=1107480 $Y=1647120
X401 1 184 189 3216 3 NOR2X1 $T=1119360 1642480 1 180 $X=1117380 $Y=1642078
X402 1 4625 365 4567 3 NOR2X1 $T=1547700 1773520 0 180 $X=1545720 $Y=1768080
X403 1 4747 421 4528 3 NOR2X1 $T=1565520 1743280 0 180 $X=1563540 $Y=1737840
X404 1 421 4692 4586 3 NOR2X1 $T=1566840 1763440 0 180 $X=1564860 $Y=1758000
X405 1 436 423 4736 3 NOR2X1 $T=1568820 1622320 0 0 $X=1568818 $Y=1621918
X406 1 452 4707 4730 3 NOR2X1 $T=1590600 1652560 0 180 $X=1588620 $Y=1647120
X407 1 453 4832 4747 3 NOR2X1 $T=1602480 1743280 0 180 $X=1600500 $Y=1737840
X408 1 459 4872 4625 3 NOR2X1 $T=1616340 1773520 0 180 $X=1614360 $Y=1768080
X409 1 4904 4706 4892 3 NOR2X1 $T=1621620 1702960 1 180 $X=1619640 $Y=1702558
X410 1 4872 4702 4905 3 NOR2X1 $T=1624260 1773520 0 180 $X=1622280 $Y=1768080
X411 1 465 4886 4949 3 NOR2X1 $T=1639440 1713040 0 0 $X=1639438 $Y=1712638
X412 1 5215 5217 5246 3 NOR2X1 $T=1727220 1692880 0 0 $X=1727218 $Y=1692478
X413 1 5319 5278 5313 3 NOR2X1 $T=1760220 1733200 0 180 $X=1758240 $Y=1727760
X414 1 5338 5305 5346 3 NOR2X1 $T=1766160 1662640 1 0 $X=1766158 $Y=1657200
X415 1 487 260 5866 3 NOR2X1 $T=1948320 1672720 0 0 $X=1948318 $Y=1672318
X416 1 5921 505 5847 3 NOR2X1 $T=1963500 1733200 1 180 $X=1961520 $Y=1732798
X417 1 5919 505 5867 3 NOR2X1 $T=1965480 1672720 0 180 $X=1963500 $Y=1667280
X418 1 5920 533 5841 3 NOR2X1 $T=1965480 1713040 1 180 $X=1963500 $Y=1712638
X419 1 614 533 5845 3 NOR2X1 $T=1970760 1723120 0 180 $X=1968780 $Y=1717680
X420 1 5929 533 5338 3 NOR2X1 $T=1980000 1662640 0 180 $X=1978020 $Y=1657200
X421 1 6181 645 6110 3 NOR2X1 $T=2062500 1753360 1 180 $X=2060520 $Y=1752958
X422 1 605 6262 6290 3 NOR2X1 $T=2108700 1753360 0 180 $X=2106720 $Y=1747920
X423 1 6366 6372 6400 3 NOR2X1 $T=2123220 1713040 1 0 $X=2123218 $Y=1707600
X424 1 6401 6459 6435 3 NOR2X1 $T=2151600 1713040 1 180 $X=2149620 $Y=1712638
X425 1 6503 6519 6533 3 NOR2X1 $T=2164140 1682800 0 0 $X=2164138 $Y=1682398
X426 1 6563 6533 6546 3 NOR2X1 $T=2172720 1672720 0 180 $X=2170740 $Y=1667280
X427 1 621 633 6637 3 NOR2X1 $T=2173380 1773520 1 0 $X=2173378 $Y=1768080
X428 1 6547 6564 6563 3 NOR2X1 $T=2175360 1682800 0 0 $X=2175358 $Y=1682398
X429 1 6621 6627 6684 3 NOR2X1 $T=2196480 1702960 0 0 $X=2196478 $Y=1702558
X430 1 6742 6684 6755 3 NOR2X1 $T=2225520 1702960 0 0 $X=2225518 $Y=1702558
X431 1 6732 6730 6742 3 NOR2X1 $T=2227500 1723120 1 180 $X=2225520 $Y=1722718
X432 1 699 6795 6844 3 NOR2X1 $T=2247300 1753360 1 0 $X=2247298 $Y=1747920
X433 1 6855 704 6858 3 NOR2X1 $T=2255220 1773520 1 0 $X=2255218 $Y=1768080
X434 1 6928 6938 713 3 NOR2X1 $T=2285580 1622320 0 0 $X=2285578 $Y=1621918
X435 1 712 7014 7028 3 NOR2X1 $T=2306700 1713040 1 0 $X=2306698 $Y=1707600
X436 1 730 728 7112 3 NOR2X1 $T=2344980 1773520 0 180 $X=2343000 $Y=1768080
X437 1 605 5936 7260 3 NOR2X1 $T=2392500 1743280 1 0 $X=2392498 $Y=1737840
X438 1 632 772 7634 3 NOR2X1 $T=2502720 1682800 0 0 $X=2502718 $Y=1682398
X439 1 798 790 800 3 NOR2X1 $T=2583240 1773520 1 180 $X=2581260 $Y=1773118
X440 1 800 801 799 3 NOR2X1 $T=2593800 1773520 0 0 $X=2593798 $Y=1773118
X441 1 7948 7925 8081 3 NOR2X1 $T=2599080 1662640 1 0 $X=2599078 $Y=1657200
X442 1 8098 7944 835 3 NOR2X1 $T=2625480 1773520 1 0 $X=2625478 $Y=1768080
X443 1896 1981 3 1 1912 NOR2X2 $T=713460 1682800 1 180 $X=710160 $Y=1682398
X444 1966 1970 3 1 1981 NOR2X2 $T=733920 1682800 0 0 $X=733918 $Y=1682398
X445 1947 1999 3 1 1983 NOR2X2 $T=739860 1723120 1 0 $X=739858 $Y=1717680
X446 2085 2080 3 1 1946 NOR2X2 $T=762960 1713040 1 0 $X=762958 $Y=1707600
X447 63 2116 3 1 2082 NOR2X2 $T=778140 1763440 1 0 $X=778138 $Y=1758000
X448 66 2144 3 1 2116 NOR2X2 $T=788040 1763440 0 180 $X=784740 $Y=1758000
X449 2494 2493 3 1 2475 NOR2X2 $T=891660 1672720 1 180 $X=888360 $Y=1672318
X450 2227 2500 3 1 2494 NOR2X2 $T=894960 1662640 1 180 $X=891660 $Y=1662238
X451 2215 2572 3 1 2493 NOR2X2 $T=895620 1692880 0 180 $X=892320 $Y=1687440
X452 3957 339 3 1 3963 NOR2X2 $T=1345740 1682800 0 0 $X=1345738 $Y=1682398
X453 3990 3963 3 1 3986 NOR2X2 $T=1351020 1672720 0 0 $X=1351018 $Y=1672318
X454 4029 4026 3 1 3990 NOR2X2 $T=1368840 1672720 1 180 $X=1365540 $Y=1672318
X455 4777 4779 3 1 4769 NOR2X2 $T=1591260 1692880 0 0 $X=1591258 $Y=1692478
X456 4702 4856 3 1 4885 NOR2X2 $T=1608420 1702960 1 0 $X=1608418 $Y=1697520
X457 5866 5867 3 1 5464 NOR2X2 $T=1950960 1672720 1 0 $X=1950958 $Y=1667280
X458 533 5933 3 1 5215 NOR2X2 $T=1960860 1692880 1 180 $X=1957560 $Y=1692478
X459 505 5936 3 1 5319 NOR2X2 $T=1969440 1733200 0 180 $X=1966140 $Y=1727760
X460 712 6945 3 1 700 NOR2X2 $T=2285580 1692880 0 180 $X=2282280 $Y=1687440
X461 5919 5929 3 1 7495 NOR2X2 $T=2471700 1723120 0 0 $X=2471698 $Y=1722718
X462 7928 7926 3 1 7980 NOR2X2 $T=2591160 1682800 1 0 $X=2591158 $Y=1677360
X463 179 185 3 1 3231 OR2XL $T=1126620 1763440 0 180 $X=1123980 $Y=1758000
X464 575 567 3 1 6621 OR2XL $T=2193180 1713040 1 0 $X=2193178 $Y=1707600
X465 561 551 3 1 6715 OR2XL $T=2204400 1682800 0 0 $X=2204398 $Y=1682398
X466 576 557 3 1 6732 OR2XL $T=2219580 1743280 1 0 $X=2219578 $Y=1737840
X467 805 8056 3 1 7989 OR2XL $T=2604360 1692880 0 180 $X=2601720 $Y=1687440
X468 1970 1966 1930 3 1 NAND2X2 $T=729960 1682800 1 0 $X=729958 $Y=1677360
X469 2006 2005 1949 3 1 NAND2X2 $T=741840 1702960 0 0 $X=741838 $Y=1702558
X470 2110 2115 2077 3 1 NAND2X2 $T=772860 1753360 1 0 $X=772858 $Y=1747920
X471 2215 2572 2516 3 1 NAND2X2 $T=903540 1692880 0 180 $X=900240 $Y=1687440
X472 2475 103 2538 3 1 NAND2X2 $T=904860 1672720 1 180 $X=901560 $Y=1672318
X473 3957 339 3954 3 1 NAND2X2 $T=1351680 1682800 0 0 $X=1351678 $Y=1682398
X474 2587 349 4117 3 1 NAND2X2 $T=1368180 1652560 0 0 $X=1368178 $Y=1652158
X475 325 362 217 3 1 NAND2X2 $T=1379400 1672720 1 180 $X=1376100 $Y=1672318
X476 4077 4065 4059 3 1 NAND2X2 $T=1382040 1642480 0 180 $X=1378740 $Y=1637040
X477 355 356 4015 3 1 NAND2X2 $T=1384020 1733200 0 0 $X=1384018 $Y=1732798
X478 332 381 3928 3 1 NAND2X2 $T=1436160 1632400 1 180 $X=1432860 $Y=1631998
X479 120 4275 382 3 1 NAND2X2 $T=1445400 1763440 1 0 $X=1445398 $Y=1758000
X480 392 122 4356 3 1 NAND2X2 $T=1462560 1753360 1 180 $X=1459260 $Y=1752958
X481 4372 4378 4370 3 1 NAND2X2 $T=1468500 1743280 0 0 $X=1468498 $Y=1742878
X482 4438 4436 393 3 1 NAND2X2 $T=1486320 1743280 0 180 $X=1483020 $Y=1737840
X483 4510 4507 4508 3 1 NAND2X2 $T=1508760 1773520 1 180 $X=1505460 $Y=1773118
X484 4581 4612 4661 3 1 NAND2X2 $T=1543740 1672720 0 180 $X=1540440 $Y=1667280
X485 4890 4872 4893 3 1 NAND2X2 $T=1619640 1733200 1 0 $X=1619638 $Y=1727760
X486 4917 4832 4888 3 1 NAND2X2 $T=1626240 1743280 1 0 $X=1626238 $Y=1737840
X487 4835 5014 5011 3 1 NAND2X2 $T=1655940 1672720 0 180 $X=1652640 $Y=1667280
X488 619 5958 618 3 1 NAND2X2 $T=1989240 1692880 1 0 $X=1989238 $Y=1687440
X489 6247 6273 651 3 1 NAND2X2 $T=2087580 1622320 1 180 $X=2084280 $Y=1621918
X490 6727 6775 694 3 1 NAND2X2 $T=2231460 1622320 1 180 $X=2228160 $Y=1621918
X491 805 8073 8043 3 1 NAND2X2 $T=2624160 1682800 0 180 $X=2620860 $Y=1677360
X492 1912 1 1949 1929 3 1931 AOI21X4 $T=726000 1702960 0 180 $X=719400 $Y=1697520
X493 1983 1 49 1948 3 46 AOI21X4 $T=735900 1723120 0 180 $X=729300 $Y=1717680
X494 2082 1 60 2077 3 1963 AOI21X4 $T=764940 1753360 0 180 $X=758340 $Y=1747920
X495 2107 1 2109 2121 3 53 AOI21X4 $T=771540 1632400 0 0 $X=771538 $Y=1631998
X496 2578 1 2476 105 3 106 AOI21X4 $T=920040 1622320 0 180 $X=913440 $Y=1616880
X497 3986 1 337 3989 3 348 AOI21X4 $T=1346400 1662640 0 0 $X=1346398 $Y=1662238
X498 350 1 4007 4020 3 4088 AOI21X4 $T=1360260 1702960 1 0 $X=1360258 $Y=1697520
X499 4077 1 4092 4096 3 4097 AOI21X4 $T=1386000 1632400 0 0 $X=1385998 $Y=1631998
X500 4397 1 123 4416 3 4349 AOI21X4 $T=1493580 1763440 0 180 $X=1486980 $Y=1758000
X501 662 1 6358 6364 3 666 AOI21X4 $T=2109360 1662640 0 0 $X=2109358 $Y=1662238
X502 696 1 6980 7015 3 6944 AOI21X4 $T=2296800 1763440 0 0 $X=2296798 $Y=1763038
X503 29 1 30 3 1765 AND2X2 $T=680460 1662640 1 180 $X=677820 $Y=1662238
X504 45 1 1945 3 43 AND2X2 $T=720060 1622320 0 180 $X=717420 $Y=1616880
X505 51 1 50 3 1978 AND2X2 $T=736560 1763440 1 180 $X=733920 $Y=1763038
X506 2027 1 1946 3 1989 AND2X2 $T=752400 1713040 0 180 $X=749760 $Y=1707600
X507 87 1 88 3 2310 AND2X2 $T=846780 1702960 1 0 $X=846778 $Y=1697520
X508 134 1 137 3 2782 AND2X2 $T=994620 1652560 1 180 $X=991980 $Y=1652158
X509 2880 1 134 3 2808 AND2X2 $T=1001220 1632400 1 180 $X=998580 $Y=1631998
X510 3150 1 3135 3 3132 AND2X2 $T=1091640 1702960 1 180 $X=1089000 $Y=1702558
X511 3231 1 3193 3 190 AND2X2 $T=1116060 1763440 0 0 $X=1116058 $Y=1763038
X512 196 1 89 3 3302 AND2X2 $T=1137840 1763440 1 0 $X=1137838 $Y=1758000
X513 210 1 268 3 3613 AND2X2 $T=1221660 1753360 0 0 $X=1221658 $Y=1752958
X514 4556 1 4559 3 4553 AND2X2 $T=1523940 1743280 1 180 $X=1521300 $Y=1742878
X515 4730 1 436 3 4658 AND2X2 $T=1567500 1642480 1 180 $X=1564860 $Y=1642078
X516 453 1 4836 3 4791 AND2X2 $T=1605120 1753360 1 180 $X=1602480 $Y=1752958
X517 456 1 380 3 4856 AND2X2 $T=1613040 1692880 1 180 $X=1610400 $Y=1692478
X518 5070 1 456 3 5038 AND2X2 $T=1686300 1692880 1 180 $X=1683660 $Y=1692478
X519 537 1 5503 3 541 AND2X2 $T=1821600 1773520 1 0 $X=1821598 $Y=1768080
X520 5529 1 5595 3 5501 AND2X2 $T=1832820 1753360 1 180 $X=1830180 $Y=1752958
X521 509 1 578 3 5614 AND2X2 $T=1863840 1682800 1 180 $X=1861200 $Y=1682398
X522 670 1 6436 3 6417 AND2X2 $T=2139060 1632400 0 180 $X=2136420 $Y=1626960
X523 700 1 6775 3 6783 AND2X2 $T=2245980 1622320 1 180 $X=2243340 $Y=1621918
X524 6775 1 6781 3 6840 AND2X2 $T=2261820 1652560 0 180 $X=2259180 $Y=1647120
X525 631 1 758 3 7550 AND2X2 $T=2509980 1702960 0 0 $X=2509978 $Y=1702558
X526 7777 1 7718 3 7719 AND2X2 $T=2532420 1642480 1 180 $X=2529780 $Y=1642078
X527 791 1 7803 3 7800 AND2X2 $T=2546940 1642480 1 180 $X=2544300 $Y=1642078
X528 7926 1 7928 3 8022 AND2X2 $T=2580600 1672720 0 0 $X=2580598 $Y=1672318
X529 8073 1 8054 3 7978 AND2X2 $T=2608980 1702960 0 180 $X=2606340 $Y=1697520
X530 8098 1 7944 3 816 AND2X2 $T=2625480 1763440 1 180 $X=2622840 $Y=1763038
X531 1912 3 1946 1 1947 NAND2X4 $T=726000 1713040 0 180 $X=721380 $Y=1707600
X532 355 3 352 1 3987 NAND2X4 $T=1376100 1723120 1 180 $X=1371480 $Y=1722718
X533 408 3 4525 1 409 NAND2X4 $T=1511400 1773520 0 0 $X=1511398 $Y=1773118
X534 4553 3 4562 1 4260 NAND2X4 $T=1521300 1733200 1 0 $X=1521298 $Y=1727760
X535 4661 3 4638 1 4522 NAND2X4 $T=1553640 1672720 1 180 $X=1549020 $Y=1672318
X536 4676 3 429 1 4686 NAND2X4 $T=1559580 1632400 1 0 $X=1559578 $Y=1626960
X537 4661 3 4715 1 4721 NAND2X4 $T=1568820 1672720 0 0 $X=1568818 $Y=1672318
X538 4888 3 4887 1 458 NAND2X4 $T=1618980 1743280 0 180 $X=1614360 $Y=1737840
X539 5261 3 352 1 5348 NAND2X4 $T=1772100 1622320 0 180 $X=1767480 $Y=1616880
X540 5261 3 362 1 5463 NAND2X4 $T=1799160 1622320 1 0 $X=1799158 $Y=1616880
X541 2054 2057 3 1 2007 OR2X2 $T=753720 1652560 0 180 $X=751080 $Y=1647120
X542 2080 2068 3 1 2006 OR2X2 $T=757680 1702960 1 180 $X=755040 $Y=1702558
X543 2116 64 3 1 2110 OR2X2 $T=774180 1763440 0 180 $X=771540 $Y=1758000
X544 2152 2118 3 1 2105 OR2X2 $T=781440 1672720 0 180 $X=778800 $Y=1667280
X545 2291 2312 3 1 2261 OR2X2 $T=836220 1743280 0 180 $X=833580 $Y=1737840
X546 2515 2533 3 1 102 OR2X2 $T=901560 1622320 0 0 $X=901558 $Y=1621918
X547 145 2898 3 1 2880 OR2X2 $T=1013760 1632400 1 180 $X=1011120 $Y=1631998
X548 156 152 3 1 2923 OR2X2 $T=1042800 1753360 1 180 $X=1040160 $Y=1752958
X549 154 153 3 1 2959 OR2X2 $T=1046760 1702960 0 180 $X=1044120 $Y=1697520
X550 3005 155 3 1 151 OR2X2 $T=1048080 1763440 1 180 $X=1045440 $Y=1763038
X551 3118 176 3 1 175 OR2X2 $T=1091640 1773520 1 180 $X=1089000 $Y=1773118
X552 184 178 3 1 3135 OR2X2 $T=1094940 1692880 1 180 $X=1092300 $Y=1692478
X553 186 179 3 1 3162 OR2X2 $T=1099560 1733200 0 180 $X=1096920 $Y=1727760
X554 178 186 3 1 3150 OR2X2 $T=1113420 1702960 1 0 $X=1113418 $Y=1697520
X555 247 227 3 1 3406 OR2X2 $T=1189320 1642480 1 180 $X=1186680 $Y=1642078
X556 229 227 3 1 3468 OR2X2 $T=1189320 1662640 0 0 $X=1189318 $Y=1662238
X557 237 227 3 1 3437 OR2X2 $T=1194600 1622320 1 180 $X=1191960 $Y=1621918
X558 239 227 3 1 3454 OR2X2 $T=1197240 1723120 0 180 $X=1194600 $Y=1717680
X559 251 242 3 1 3481 OR2X2 $T=1201200 1642480 0 180 $X=1198560 $Y=1637040
X560 258 242 3 1 3438 OR2X2 $T=1202520 1632400 0 180 $X=1199880 $Y=1626960
X561 260 242 3 1 3471 OR2X2 $T=1213080 1682800 1 180 $X=1210440 $Y=1682398
X562 272 242 3 1 3462 OR2X2 $T=1230900 1723120 1 180 $X=1228260 $Y=1722718
X563 2743 344 3 1 4007 OR2X2 $T=1345080 1702960 1 0 $X=1345078 $Y=1697520
X564 4241 375 3 1 4228 OR2X2 $T=1432860 1652560 1 180 $X=1430220 $Y=1652158
X565 4767 4625 3 1 4773 OR2X2 $T=1589280 1763440 0 0 $X=1589278 $Y=1763038
X566 450 441 3 1 4774 OR2X2 $T=1590600 1642480 1 0 $X=1590598 $Y=1637040
X567 456 380 3 1 4886 OR2X2 $T=1610400 1713040 0 0 $X=1610398 $Y=1712638
X568 582 595 3 1 5767 OR2X2 $T=1914660 1652560 1 0 $X=1914658 $Y=1647120
X569 341 487 3 1 5768 OR2X2 $T=1924560 1743280 1 180 $X=1921920 $Y=1742878
X570 533 605 3 1 5758 OR2X2 $T=1948980 1753360 1 180 $X=1946340 $Y=1752958
X571 533 610 3 1 609 OR2X2 $T=1963500 1622320 0 180 $X=1960860 $Y=1616880
X572 505 5900 3 1 5309 OR2X2 $T=1968780 1682800 1 180 $X=1966140 $Y=1682398
X573 6259 6218 3 1 6247 OR2X2 $T=2084280 1642480 0 180 $X=2081640 $Y=1637040
X574 655 6246 3 1 6245 OR2X2 $T=2086260 1723120 1 180 $X=2083620 $Y=1722718
X575 653 6257 3 1 6224 OR2X2 $T=2088900 1692880 1 180 $X=2086260 $Y=1692478
X576 658 6291 3 1 6268 OR2X2 $T=2099460 1622320 1 180 $X=2096820 $Y=1621918
X577 661 6341 3 1 6250 OR2X2 $T=2110020 1642480 1 180 $X=2107380 $Y=1642078
X578 664 667 3 1 6358 OR2X2 $T=2128500 1672720 0 180 $X=2125860 $Y=1667280
X579 5921 6342 3 1 6366 OR2X2 $T=2131140 1723120 0 180 $X=2128500 $Y=1717680
X580 678 673 3 1 670 OR2X2 $T=2145000 1632400 0 180 $X=2142360 $Y=1626960
X581 6679 6608 3 1 6567 OR2X2 $T=2201760 1662640 0 180 $X=2199120 $Y=1657200
X582 6785 6772 3 1 6857 OR2X2 $T=2238060 1682800 1 0 $X=2238058 $Y=1677360
X583 6891 6874 3 1 6775 OR2X2 $T=2264460 1652560 0 180 $X=2261820 $Y=1647120
X584 6909 6907 3 1 6932 OR2X2 $T=2275020 1702960 0 0 $X=2275018 $Y=1702558
X585 7040 7029 3 1 720 OR2X2 $T=2310000 1622320 0 180 $X=2307360 $Y=1616880
X586 7086 7045 3 1 6959 OR2X2 $T=2327820 1692880 0 180 $X=2325180 $Y=1687440
X587 8095 7963 3 1 8073 OR2X2 $T=2624160 1702960 1 0 $X=2624158 $Y=1697520
X588 2247 3 1 2275 2273 NAND2XL $T=829620 1652560 1 180 $X=827640 $Y=1652158
X589 2275 3 1 71 2272 NAND2XL $T=835560 1652560 1 0 $X=835558 $Y=1647120
X590 2310 3 1 85 2393 NAND2XL $T=854700 1672720 0 0 $X=854698 $Y=1672318
X591 2310 3 1 86 2392 NAND2XL $T=856020 1662640 0 0 $X=856018 $Y=1662238
X592 86 3 1 85 2391 NAND2XL $T=865920 1662640 0 180 $X=863940 $Y=1657200
X593 2227 3 1 2500 2510 NAND2XL $T=892980 1652560 0 0 $X=892978 $Y=1652158
X594 2983 3 1 2959 2947 NAND2XL $T=1030920 1702960 0 180 $X=1028940 $Y=1697520
X595 178 3 1 184 3187 NAND2XL $T=1100880 1692880 0 0 $X=1100878 $Y=1692478
X596 185 3 1 183 3152 NAND2XL $T=1102860 1642480 0 180 $X=1100880 $Y=1637040
X597 4117 3 1 4065 4170 NAND2XL $T=1403820 1642480 1 0 $X=1403818 $Y=1637040
X598 422 3 1 5020 5036 NAND2XL $T=1657920 1763440 1 0 $X=1657918 $Y=1758000
X599 6181 3 1 645 6112 NAND2XL $T=2065140 1753360 1 180 $X=2063160 $Y=1752958
X600 6212 3 1 6224 6221 NAND2XL $T=2076360 1702960 0 0 $X=2076358 $Y=1702558
X601 6325 3 1 6268 6292 NAND2XL $T=2102100 1642480 0 180 $X=2100120 $Y=1637040
X602 6608 3 1 6679 6617 NAND2XL $T=2204400 1662640 1 0 $X=2204398 $Y=1657200
X603 6621 3 1 6627 6705 NAND2XL $T=2207040 1702960 0 0 $X=2207038 $Y=1702558
X604 549 3 1 6715 6729 NAND2XL $T=2218920 1682800 1 0 $X=2218918 $Y=1677360
X605 6724 3 1 6727 6739 NAND2XL $T=2220240 1632400 1 0 $X=2220238 $Y=1626960
X606 6732 3 1 6730 6712 NAND2XL $T=2222220 1723120 0 180 $X=2220240 $Y=1717680
X607 699 3 1 6795 6842 NAND2XL $T=2240040 1753360 1 0 $X=2240038 $Y=1747920
X608 6755 3 1 6799 6785 NAND2XL $T=2241360 1702960 0 0 $X=2241358 $Y=1702558
X609 7065 3 1 6959 7044 NAND2XL $T=2327820 1702960 0 180 $X=2325840 $Y=1697520
X610 2515 2578 3 1 INVX4 $T=914760 1632400 0 0 $X=914758 $Y=1631998
X611 231 215 3 1 INVX4 $T=1189980 1632400 0 0 $X=1189978 $Y=1631998
X612 4524 4552 3 1 INVX4 $T=1519980 1702960 1 0 $X=1519978 $Y=1697520
X613 4572 4849 3 1 INVX4 $T=1618320 1682800 0 0 $X=1618318 $Y=1682398
X614 4706 4917 3 1 INVX4 $T=1628880 1723120 0 180 $X=1626240 $Y=1717680
X615 484 5261 3 1 INVX4 $T=1712700 1622320 1 0 $X=1712698 $Y=1616880
X616 5715 567 3 1 INVX4 $T=1893540 1632400 1 180 $X=1890900 $Y=1631998
X617 582 591 3 1 INVX4 $T=1910040 1763440 0 0 $X=1910038 $Y=1763038
X618 6096 5919 3 1 INVX4 $T=2044680 1672720 1 0 $X=2044678 $Y=1667280
X619 5973 6166 3 1 INVX4 $T=2051280 1702960 0 0 $X=2051278 $Y=1702558
X620 668 602 3 1 INVX4 $T=2167440 1743280 1 180 $X=2164800 $Y=1742878
X621 621 614 3 1 INVX4 $T=2176020 1723120 1 180 $X=2173380 $Y=1722718
X622 623 5921 3 1 INVX4 $T=2361480 1723120 0 180 $X=2358840 $Y=1717680
X623 632 610 3 1 INVX4 $T=2429460 1622320 1 0 $X=2429458 $Y=1616880
X624 1946 1964 1 1949 1982 3 AOI21X1 $T=728640 1713040 1 0 $X=728638 $Y=1707600
X625 50 51 1 48 1928 3 AOI21X1 $T=734580 1773520 1 0 $X=734578 $Y=1768080
X626 65 67 1 2150 2156 3 AOI21X1 $T=788040 1773520 0 0 $X=788038 $Y=1773118
X627 2245 70 1 2258 2244 3 AOI21X1 $T=813780 1763440 1 0 $X=813778 $Y=1758000
X628 2258 2261 1 2262 2228 3 AOI21X1 $T=820380 1743280 0 180 $X=817740 $Y=1737840
X629 94 2542 1 2543 2550 3 AOI21X1 $T=904860 1702960 1 0 $X=904858 $Y=1697520
X630 83 2509 1 107 2591 3 AOI21X1 $T=915420 1763440 0 0 $X=915418 $Y=1763038
X631 2604 2477 1 2606 2608 3 AOI21X1 $T=922680 1733200 0 0 $X=922678 $Y=1732798
X632 134 2809 1 2805 2801 3 AOI21X1 $T=991980 1642480 1 180 $X=989340 $Y=1642078
X633 2805 2880 1 2883 2804 3 AOI21X1 $T=1006500 1642480 1 0 $X=1006498 $Y=1637040
X634 2925 2923 1 2922 2919 3 AOI21X1 $T=1019040 1763440 0 180 $X=1016400 $Y=1758000
X635 151 150 1 2925 146 3 AOI21X1 $T=1034880 1773520 1 180 $X=1032240 $Y=1773118
X636 3214 3135 1 3203 3165 3 AOI21X1 $T=1108140 1702960 1 180 $X=1105500 $Y=1702558
X637 3150 3161 1 3214 3189 3 AOI21X1 $T=1109460 1713040 0 180 $X=1106820 $Y=1707600
X638 274 273 1 3613 271 3 AOI21X1 $T=1232220 1753360 0 180 $X=1229580 $Y=1747920
X639 4065 4131 1 4092 361 3 AOI21X1 $T=1397220 1632400 0 0 $X=1397218 $Y=1631998
X640 373 4253 1 372 378 3 AOI21X1 $T=1438140 1662640 0 180 $X=1435500 $Y=1657200
X641 4419 4512 1 4514 4507 3 AOI21X1 $T=1509420 1723120 1 0 $X=1509418 $Y=1717680
X642 4437 4512 1 4514 4513 3 AOI21X1 $T=1510080 1733200 1 0 $X=1510078 $Y=1727760
X643 441 4736 1 4738 4729 3 AOI21X1 $T=1577400 1642480 1 0 $X=1577398 $Y=1637040
X644 4791 4773 1 421 4770 3 AOI21X1 $T=1592580 1753360 1 180 $X=1589940 $Y=1752958
X645 5548 5556 1 5561 568 3 AOI21X1 $T=1846020 1773520 1 0 $X=1846018 $Y=1768080
X646 525 563 1 5566 5548 3 AOI21X1 $T=1849980 1723120 0 180 $X=1847340 $Y=1717680
X647 6224 6215 1 6219 6218 3 AOI21X1 $T=2077680 1692880 1 180 $X=2075040 $Y=1692478
X648 6250 6256 1 6261 6293 3 AOI21X1 $T=2087580 1652560 0 0 $X=2087578 $Y=1652158
X649 6261 6268 1 6269 6273 3 AOI21X1 $T=2090220 1632400 1 0 $X=2090218 $Y=1626960
X650 670 6392 1 6389 6391 3 AOI21X1 $T=2125860 1622320 1 180 $X=2123220 $Y=1621918
X651 6326 6439 1 6441 6521 3 AOI21X1 $T=2138400 1692880 1 0 $X=2138398 $Y=1687440
X652 6471 6470 1 6468 6469 3 AOI21X1 $T=2148960 1662640 1 180 $X=2146320 $Y=1662238
X653 6567 6549 1 6593 6576 3 AOI21X1 $T=2183280 1652560 0 0 $X=2183278 $Y=1652158
X654 6767 6755 1 6711 6764 3 AOI21X1 $T=2232780 1702960 1 180 $X=2230140 $Y=1702558
X655 766 767 1 5936 7579 3 AOI21X1 $T=2490840 1642480 1 0 $X=2490838 $Y=1637040
X656 42 1928 3 41 1 1884 OAI21X2 $T=710820 1773520 0 180 $X=705540 $Y=1768080
X657 2243 69 3 2228 1 2109 OAI21X2 $T=810480 1733200 1 180 $X=805200 $Y=1732798
X658 2493 2614 3 2516 1 2577 OAI21X2 $T=920040 1682800 0 180 $X=914760 $Y=1677360
X659 3954 3990 3 4010 1 3989 OAI21X2 $T=1356960 1672720 1 0 $X=1356958 $Y=1667280
X660 4781 4857 3 4770 1 4743 OAI21X2 $T=1595880 1733200 1 180 $X=1590600 $Y=1732798
X661 4857 4905 3 459 1 461 OAI21X2 $T=1624920 1773520 1 180 $X=1619640 $Y=1773118
X662 5921 614 3 6977 1 7023 OAI21X2 $T=2302740 1733200 0 180 $X=2297460 $Y=1727760
X663 40 1884 1895 3 1 XNOR2X4 $T=702240 1753360 0 0 $X=702238 $Y=1752958
X664 1917 1961 57 3 1 XNOR2X4 $T=726000 1652560 0 0 $X=725998 $Y=1652158
X665 6947 6944 710 3 1 XNOR2X4 $T=2290860 1773520 0 180 $X=2279640 $Y=1768080
X666 1963 3 1947 1931 1 1948 OAI21X4 $T=725340 1713040 1 180 $X=718080 $Y=1712638
X667 4059 3 4088 4097 1 357 OAI21X4 $T=1385340 1642480 0 0 $X=1385338 $Y=1642078
X668 4327 3 4323 157 1 4321 OAI21X4 $T=1454640 1753360 1 180 $X=1447380 $Y=1752958
X669 4397 3 4387 130 1 4340 OAI21X4 $T=1473120 1743280 0 0 $X=1473118 $Y=1742878
X670 399 3 398 387 1 4460 OAI21X4 $T=1497540 1652560 0 180 $X=1490280 $Y=1647120
X671 399 3 398 4500 1 4471 OAI21X4 $T=1500840 1672720 1 0 $X=1500838 $Y=1667280
X672 6945 3 714 6971 1 701 OAI21X4 $T=2290860 1692880 1 0 $X=2290858 $Y=1687440
X673 2643 3 30 1 CLKBUFX8 $T=937860 1763440 0 180 $X=933240 $Y=1758000
X674 2715 3 119 1 CLKBUFX8 $T=961620 1622320 1 0 $X=961618 $Y=1616880
X675 2803 3 37 1 CLKBUFX8 $T=993960 1743280 1 0 $X=993958 $Y=1737840
X676 2989 3 27 1 CLKBUFX8 $T=1046100 1642480 0 0 $X=1046098 $Y=1642078
X677 3077 3 29 1 CLKBUFX8 $T=1077120 1652560 1 0 $X=1077118 $Y=1647120
X678 3075 3 28 1 CLKBUFX8 $T=1077780 1692880 1 0 $X=1077778 $Y=1687440
X679 3369 3 104 1 CLKBUFX8 $T=1160280 1702960 0 180 $X=1155660 $Y=1697520
X680 3639 3 278 1 CLKBUFX8 $T=1238160 1642480 1 180 $X=1233540 $Y=1642078
X681 3733 3 184 1 CLKBUFX8 $T=1270500 1662640 1 180 $X=1265880 $Y=1662238
X682 5261 3 514 1 CLKBUFX8 $T=1774740 1622320 1 0 $X=1774738 $Y=1616880
X683 5381 3 5393 1 CLKBUFX8 $T=1782000 1682800 0 0 $X=1781998 $Y=1682398
X684 5456 3 533 1 CLKBUFX8 $T=1801800 1622320 0 0 $X=1801798 $Y=1621918
X685 5348 3 538 1 CLKBUFX8 $T=1816320 1622320 1 0 $X=1816318 $Y=1616880
X686 5463 3 550 1 CLKBUFX8 $T=1820940 1622320 1 0 $X=1820938 $Y=1616880
X687 6059 3 633 1 CLKBUFX8 $T=2022240 1723120 0 0 $X=2022238 $Y=1722718
X688 6046 3 623 1 CLKBUFX8 $T=2026200 1733200 0 0 $X=2026198 $Y=1732798
X689 1953 1960 1 3 1966 XOR2X2 $T=726000 1743280 0 0 $X=725998 $Y=1742878
X690 1962 1969 1 3 52 XOR2X2 $T=729300 1662640 0 0 $X=729298 $Y=1662238
X691 2104 2139 1 3 2154 XOR2X2 $T=783420 1692880 1 0 $X=783418 $Y=1687440
X692 2168 2156 1 3 2215 XOR2X2 $T=793320 1743280 1 0 $X=793318 $Y=1737840
X693 2590 2614 1 3 2743 XOR2X2 $T=924660 1692880 1 0 $X=924658 $Y=1687440
X694 6399 6391 1 3 368 XOR2X2 $T=2127180 1622320 0 180 $X=2120580 $Y=1616880
X695 6417 6392 1 3 4029 XOR2X2 $T=2131800 1632400 0 180 $X=2125200 $Y=1626960
X696 7222 7221 1 3 730 XOR2X2 $T=2383260 1702960 1 180 $X=2376660 $Y=1702558
X697 7989 7978 1 3 6909 XOR2X2 $T=2599080 1702960 0 180 $X=2592480 $Y=1697520
X698 8026 8023 1 3 6728 XOR2X2 $T=2603700 1652560 0 180 $X=2597100 $Y=1647120
X699 88 3 98 1 INVX2 $T=914100 1753360 0 180 $X=912120 $Y=1747920
X700 2781 3 2809 1 INVX2 $T=985380 1662640 1 0 $X=985378 $Y=1657200
X701 222 3 347 1 INVX2 $T=1378080 1662640 1 0 $X=1378078 $Y=1657200
X702 287 3 282 1 INVX2 $T=1395240 1733200 1 0 $X=1395238 $Y=1727760
X703 300 3 307 1 INVX2 $T=1401180 1713040 1 0 $X=1401178 $Y=1707600
X704 220 3 235 1 INVX2 $T=1411740 1723120 0 0 $X=1411738 $Y=1722718
X705 234 3 233 1 INVX2 $T=1440780 1702960 1 0 $X=1440778 $Y=1697520
X706 221 3 257 1 INVX2 $T=1444740 1632400 1 0 $X=1444738 $Y=1626960
X707 236 3 261 1 INVX2 $T=1482360 1642480 0 0 $X=1482358 $Y=1642078
X708 213 3 203 1 INVX2 $T=1495560 1692880 0 0 $X=1495558 $Y=1692478
X709 230 3 223 1 INVX2 $T=1509420 1682800 1 0 $X=1509418 $Y=1677360
X710 4540 3 4477 1 INVX2 $T=1519320 1743280 1 0 $X=1519318 $Y=1737840
X711 415 3 4716 1 INVX2 $T=1571460 1713040 0 0 $X=1571458 $Y=1712638
X712 4893 3 4895 1 INVX2 $T=1618980 1743280 1 0 $X=1618978 $Y=1737840
X713 666 3 6392 1 INVX2 $T=2131140 1622320 0 0 $X=2131138 $Y=1621918
X714 631 3 7262 1 INVX2 $T=2436720 1652560 1 180 $X=2434740 $Y=1652158
X715 90 1 3 2410 INVXL $T=852720 1713040 0 0 $X=852718 $Y=1712638
X716 2900 1 3 2865 INVXL $T=1003200 1713040 1 180 $X=1001880 $Y=1712638
X717 34 1 3 3356 INVXL $T=1143120 1753360 1 0 $X=1143118 $Y=1747920
X718 97 1 3 3516 INVXL $T=1200540 1743280 1 0 $X=1200538 $Y=1737840
X719 337 1 3 3894 INVXL $T=1323300 1682800 0 0 $X=1323298 $Y=1682398
X720 375 1 3 4253 INVXL $T=1438140 1672720 1 0 $X=1438138 $Y=1667280
X721 123 1 3 4378 INVXL $T=1474440 1753360 0 180 $X=1473120 $Y=1747920
X722 4918 1 3 4884 INVXL $T=1618980 1642480 0 180 $X=1617660 $Y=1637040
X723 594 1 3 5500 INVXL $T=1884300 1652560 0 180 $X=1882980 $Y=1647120
X724 5919 1 3 6055 INVXL $T=2049300 1642480 1 180 $X=2047980 $Y=1642078
X725 6505 1 3 6468 INVXL $T=2153580 1662640 1 180 $X=2152260 $Y=1662238
X726 6533 1 3 6471 INVXL $T=2156220 1672720 0 180 $X=2154900 $Y=1667280
X727 6742 1 3 6747 INVXL $T=2225520 1723120 1 0 $X=2225518 $Y=1717680
X728 6767 1 3 6870 INVXL $T=2250600 1723120 1 0 $X=2250598 $Y=1717680
X729 122 4415 4403 1 4400 4322 3 AOI31X1 $T=1481700 1733200 0 180 $X=1478400 $Y=1727760
X730 1927 45 1 3 1894 XNOR2X2 $T=720060 1642480 0 180 $X=712800 $Y=1637040
X731 2571 2577 1 3 2587 XNOR2X2 $T=913440 1652560 0 0 $X=913438 $Y=1652158
X732 2585 2578 1 3 2620 XNOR2X2 $T=920700 1622320 0 0 $X=920698 $Y=1621918
X733 662 6354 1 3 3957 XNOR2X2 $T=2112000 1682800 1 180 $X=2104740 $Y=1682398
X734 6840 6841 1 3 6032 XNOR2X2 $T=2251920 1652560 0 180 $X=2244660 $Y=1647120
X735 621 6166 1 3 7372 XNOR2X2 $T=2434740 1672720 1 0 $X=2434738 $Y=1667280
X736 2106 2094 3 1 2114 XOR2X1 $T=770880 1692880 1 0 $X=770878 $Y=1687440
X737 2246 2244 3 1 2144 XOR2X1 $T=813120 1753360 1 180 $X=807840 $Y=1752958
X738 2249 2247 3 1 2217 XOR2X1 $T=815100 1662640 1 180 $X=809820 $Y=1662238
X739 71 2275 3 1 2249 XOR2X1 $T=823020 1662640 0 180 $X=817740 $Y=1657200
X740 2311 2310 3 1 2275 XOR2X1 $T=836220 1662640 1 180 $X=830940 $Y=1662238
X741 85 86 3 1 2311 XOR2X1 $T=846780 1662640 1 180 $X=841500 $Y=1662238
X742 88 87 3 1 2322 XOR2X1 $T=859980 1723120 1 180 $X=854700 $Y=1722718
X743 2815 2801 3 1 2572 XOR2X1 $T=997260 1662640 1 180 $X=991980 $Y=1662238
X744 2915 2900 3 1 141 XOR2X1 $T=1017060 1743280 0 180 $X=1011780 $Y=1737840
X745 167 168 3 1 2898 XOR2X1 $T=1069200 1632400 0 180 $X=1063920 $Y=1626960
X746 3192 3189 3 1 180 XOR2X1 $T=1105500 1713040 1 180 $X=1100220 $Y=1712638
X747 3193 3190 3 1 181 XOR2X1 $T=1105500 1763440 1 180 $X=1100220 $Y=1763038
X748 3211 3197 3 1 3118 XOR2X1 $T=1108140 1672720 1 180 $X=1102860 $Y=1672318
X749 3898 3894 3 1 335 XOR2X1 $T=1325280 1672720 1 180 $X=1320000 $Y=1672318
X750 372 4228 3 1 370 XOR2X1 $T=1427580 1652560 1 180 $X=1422300 $Y=1652158
X751 4241 375 3 1 379 XOR2X1 $T=1434840 1652560 0 0 $X=1434838 $Y=1652158
X752 456 380 3 1 4946 XOR2X1 $T=1634160 1692880 0 0 $X=1634158 $Y=1692478
X753 639 6098 3 1 637 XOR2X1 $T=2040720 1763440 1 180 $X=2035440 $Y=1763038
X754 6183 6182 3 1 644 XOR2X1 $T=2065800 1743280 0 180 $X=2060520 $Y=1737840
X755 6248 6256 3 1 650 XOR2X1 $T=2089560 1662640 1 180 $X=2084280 $Y=1662238
X756 6292 6293 3 1 659 XOR2X1 $T=2097480 1662640 1 0 $X=2097478 $Y=1657200
X757 6418 6409 3 1 6323 XOR2X1 $T=2131800 1702960 1 180 $X=2126520 $Y=1702558
X758 6479 6469 3 1 6410 XOR2X1 $T=2151600 1652560 1 180 $X=2146320 $Y=1652158
X759 6552 6551 3 1 6544 XOR2X1 $T=2172720 1642480 0 180 $X=2167440 $Y=1637040
X760 6622 6619 3 1 687 XOR2X1 $T=2196480 1773520 1 180 $X=2191200 $Y=1773118
X761 6901 695 3 1 6907 XOR2X1 $T=2269740 1733200 1 0 $X=2269738 $Y=1727760
X762 6888 6908 3 1 7045 XOR2X1 $T=2275020 1753360 1 0 $X=2275018 $Y=1747920
X763 7187 718 3 1 7222 XOR2X1 $T=2376660 1692880 0 0 $X=2376658 $Y=1692478
X764 7013 6507 3 1 742 XOR2X1 $T=2376660 1753360 0 0 $X=2376658 $Y=1752958
X765 7248 7250 3 1 7221 XOR2X1 $T=2397780 1692880 0 180 $X=2392500 $Y=1687440
X766 7332 7331 3 1 7327 XOR2X1 $T=2416260 1753360 1 180 $X=2410980 $Y=1752958
X767 7347 7329 3 1 7332 XOR2X1 $T=2418900 1753360 0 180 $X=2413620 $Y=1747920
X768 7372 5929 3 1 7248 XOR2X1 $T=2426820 1672720 1 180 $X=2421540 $Y=1672318
X769 7191 7395 3 1 757 XOR2X1 $T=2439360 1743280 0 0 $X=2439358 $Y=1742878
X770 7465 632 3 1 755 XOR2X1 $T=2452560 1753360 1 180 $X=2447280 $Y=1752958
X771 7333 7416 3 1 7491 XOR2X1 $T=2449920 1692880 1 0 $X=2449918 $Y=1687440
X772 7492 7494 3 1 7508 XOR2X1 $T=2460480 1692880 1 0 $X=2460478 $Y=1687440
X773 7372 626 3 1 7479 XOR2X1 $T=2463120 1672720 1 0 $X=2463118 $Y=1667280
X774 7509 6342 3 1 760 XOR2X1 $T=2468400 1743280 1 180 $X=2463120 $Y=1742878
X775 7491 7508 3 1 764 XOR2X1 $T=2468400 1692880 1 0 $X=2468398 $Y=1687440
X776 614 7637 3 1 770 XOR2X1 $T=2504700 1763440 0 180 $X=2499420 $Y=1758000
X777 7578 772 3 1 7635 XOR2X1 $T=2500740 1622320 1 0 $X=2500738 $Y=1616880
X778 7660 631 3 1 7721 XOR2X1 $T=2508660 1763440 0 0 $X=2508658 $Y=1763038
X779 7701 623 3 1 779 XOR2X1 $T=2520540 1682800 0 180 $X=2515260 $Y=1677360
X780 7746 632 3 1 7804 XOR2X1 $T=2528460 1672720 0 0 $X=2528458 $Y=1672318
X781 7812 756 3 1 7836 XOR2X1 $T=2544300 1652560 0 0 $X=2544298 $Y=1652158
X782 634 613 3 1 7864 XOR2X1 $T=2559480 1632400 0 0 $X=2559478 $Y=1631998
X783 7897 7701 3 1 7926 XOR2X1 $T=2567400 1672720 1 0 $X=2567398 $Y=1667280
X784 7931 7929 3 1 798 XOR2X1 $T=2580600 1763440 1 0 $X=2580598 $Y=1758000
X785 797 7644 3 1 7929 XOR2X1 $T=2585880 1743280 0 180 $X=2580600 $Y=1737840
X786 8086 821 3 1 834 XOR2X1 $T=2623500 1723120 1 0 $X=2623498 $Y=1717680
X787 8059 820 3 1 821 XOR2X1 $T=2625480 1713040 0 0 $X=2625478 $Y=1712638
X788 2137 1 2140 2164 3 NOR2BX1 $T=792660 1713040 0 0 $X=792658 $Y=1712638
X789 389 1 4418 4416 3 NOR2BX1 $T=1485000 1763440 0 180 $X=1482360 $Y=1758000
X790 387 1 406 4500 3 NOR2BX1 $T=1506120 1662640 0 180 $X=1503480 $Y=1657200
X791 457 1 4755 4851 3 NOR2BX1 $T=1613040 1753360 0 180 $X=1610400 $Y=1747920
X792 460 1 448 4918 3 NOR2BX1 $T=1626240 1632400 0 0 $X=1626238 $Y=1631998
X793 486 1 487 5217 3 NOR2BX1 $T=1727880 1713040 1 0 $X=1727878 $Y=1707600
X794 473 1 487 5305 3 NOR2BX1 $T=1735800 1662640 1 0 $X=1735798 $Y=1657200
X795 5280 1 487 5278 3 NOR2BX1 $T=1750320 1733200 0 180 $X=1747680 $Y=1727760
X796 6442 1 6435 6418 3 NOR2BX1 $T=2138400 1702960 1 180 $X=2135760 $Y=1702558
X797 6842 1 6844 6888 3 NOR2BX1 $T=2253900 1753360 1 0 $X=2253898 $Y=1747920
X798 7527 1 7550 7511 3 NOR2BX1 $T=2480280 1702960 0 0 $X=2480278 $Y=1702558
X799 8020 1 7943 8026 3 NOR2BX1 $T=2599080 1642480 0 0 $X=2599078 $Y=1642078
X800 31 27 1765 21 1 3 2 ADDFX2 $T=674520 1632400 0 180 $X=660660 $Y=1626960
X801 34 33 28 26 1 3 22 ADDFX2 $T=681120 1702960 0 180 $X=667260 $Y=1697520
X802 2304 2322 2307 2226 1 3 2113 ADDFX2 $T=842160 1672720 1 180 $X=828300 $Y=1672318
X803 87 84 80 76 1 3 2290 ADDFX2 $T=842820 1632400 1 180 $X=828960 $Y=1631998
X804 2336 2290 81 2014 1 3 2171 ADDFX2 $T=842820 1642480 0 180 $X=828960 $Y=1637040
X805 2310 83 2301 2133 1 3 2291 ADDFX2 $T=842820 1713040 0 180 $X=828960 $Y=1707600
X806 89 85 82 2304 1 3 2301 ADDFX2 $T=843480 1682800 1 180 $X=829620 $Y=1682398
X807 85 86 83 78 1 3 74 ADDFX2 $T=844140 1622320 0 180 $X=830280 $Y=1616880
X808 83 91 2382 2347 1 3 2302 ADDFX2 $T=858660 1753360 0 180 $X=844800 $Y=1747920
X809 2410 84 2322 2312 1 3 2352 ADDFX2 $T=861300 1733200 1 180 $X=847440 $Y=1732798
X810 95 94 92 2247 1 3 2307 ADDFX2 $T=865920 1642480 0 180 $X=852060 $Y=1637040
X811 84 95 2422 75 1 3 93 ADDFX2 $T=876480 1773520 1 180 $X=862620 $Y=1773118
X812 5053 5042 471 469 1 3 468 ADDFX2 $T=1669800 1652560 1 180 $X=1655940 $Y=1652158
X813 5920 668 608 6401 1 3 6372 ADDFX2 $T=2137740 1733200 0 180 $X=2123880 $Y=1727760
X814 5936 621 5814 6503 1 3 6459 ADDFX2 $T=2164140 1723120 1 180 $X=2150280 $Y=1722718
X815 5933 623 602 6547 1 3 6519 ADDFX2 $T=2158200 1692880 1 0 $X=2158198 $Y=1687440
X816 5921 5929 6935 6928 1 3 6679 ADDFX2 $T=2292840 1662640 1 180 $X=2278980 $Y=1662238
X817 6979 5900 7024 7029 1 3 6938 ADDFX2 $T=2298120 1652560 0 0 $X=2298118 $Y=1652158
X818 610 6342 5936 723 1 3 7062 ADDFX2 $T=2335080 1642480 0 180 $X=2321220 $Y=1637040
X819 7066 7085 7062 724 1 3 7040 ADDFX2 $T=2336400 1632400 0 180 $X=2322540 $Y=1626960
X820 727 6507 5920 7066 1 3 7024 ADDFX2 $T=2337060 1652560 1 180 $X=2323200 $Y=1652158
X821 7171 6507 6166 731 1 3 729 ADDFX2 $T=2361480 1662640 0 180 $X=2347620 $Y=1657200
X822 6342 631 5919 734 1 3 732 ADDFX2 $T=2363460 1632400 1 180 $X=2349600 $Y=1631998
X823 623 6507 5929 7152 1 3 736 ADDFX2 $T=2368080 1652560 0 180 $X=2354220 $Y=1647120
X824 739 7152 7258 743 1 3 745 ADDFX2 $T=2385240 1622320 0 0 $X=2385238 $Y=1621918
X825 633 6342 7262 744 1 3 7258 ADDFX2 $T=2408340 1642480 1 180 $X=2394480 $Y=1642078
X826 55 51 3 1 2055 XNOR2X1 $T=745140 1773520 1 0 $X=745138 $Y=1768080
X827 2084 2083 3 1 2059 XNOR2X1 $T=764940 1682800 0 180 $X=759660 $Y=1677360
X828 131 129 3 1 2500 XNOR2X1 $T=985380 1632400 1 180 $X=980100 $Y=1631998
X829 2782 2781 3 1 128 XNOR2X1 $T=985380 1682800 1 180 $X=980100 $Y=1682398
X830 2862 2830 3 1 135 XNOR2X1 $T=1000560 1713040 0 180 $X=995280 $Y=1707600
X831 2947 2946 3 1 140 XNOR2X1 $T=1026960 1723120 1 180 $X=1021680 $Y=1722718
X832 3122 3120 3 1 3005 XNOR2X1 $T=1087020 1672720 0 180 $X=1081740 $Y=1667280
X833 3225 3161 3 1 188 XNOR2X1 $T=1110780 1733200 1 0 $X=1110778 $Y=1727760
X834 3948 3936 3 1 330 XNOR2X1 $T=1343760 1662640 0 180 $X=1338480 $Y=1657200
X835 4030 350 3 1 4026 XNOR2X1 $T=1369500 1702960 0 0 $X=1369498 $Y=1702558
X836 4170 4131 3 1 367 XNOR2X1 $T=1403820 1632400 1 0 $X=1403818 $Y=1626960
X837 469 477 3 1 475 XNOR2X1 $T=1686300 1642480 0 180 $X=1681020 $Y=1637040
X838 587 589 3 1 5042 XNOR2X1 $T=1906080 1652560 1 180 $X=1900800 $Y=1652158
X839 6215 6221 3 1 647 XNOR2X1 $T=2077680 1723120 0 180 $X=2072400 $Y=1717680
X840 6342 5921 3 1 6262 XNOR2X1 $T=2110020 1733200 1 180 $X=2104740 $Y=1732798
X841 6478 6470 3 1 6452 XNOR2X1 $T=2151600 1652560 0 180 $X=2146320 $Y=1647120
X842 6637 6507 3 1 6619 XNOR2X1 $T=2199120 1763440 1 180 $X=2193840 $Y=1763038
X843 567 575 3 1 6730 XNOR2X1 $T=2209020 1723120 0 0 $X=2209018 $Y=1722718
X844 6754 6766 3 1 697 XNOR2X1 $T=2230140 1662640 0 0 $X=2230138 $Y=1662238
X845 6748 6871 3 1 6874 XNOR2X1 $T=2259180 1713040 1 0 $X=2259178 $Y=1707600
X846 623 6166 3 1 6976 XNOR2X1 $T=2317920 1723120 1 180 $X=2312640 $Y=1722718
X847 633 5814 3 1 7013 XNOR2X1 $T=2313960 1733200 0 0 $X=2313958 $Y=1732798
X848 6976 5920 3 1 7049 XNOR2X1 $T=2313960 1743280 1 0 $X=2313958 $Y=1737840
X849 726 7070 3 1 722 XNOR2X1 $T=2331120 1773520 1 180 $X=2325840 $Y=1773118
X850 7185 5936 3 1 7160 XNOR2X1 $T=2368740 1733200 1 180 $X=2363460 $Y=1732798
X851 633 5919 3 1 7185 XNOR2X1 $T=2376660 1723120 1 180 $X=2371380 $Y=1722718
X852 7262 6507 3 1 7301 XNOR2X1 $T=2396460 1733200 1 0 $X=2396458 $Y=1727760
X853 7333 718 3 1 7329 XNOR2X1 $T=2413620 1702960 1 0 $X=2413618 $Y=1697520
X854 668 5936 3 1 7191 XNOR2X1 $T=2431440 1743280 0 180 $X=2426160 $Y=1737840
X855 623 5919 3 1 7333 XNOR2X1 $T=2428800 1692880 1 0 $X=2428798 $Y=1687440
X856 5929 7313 3 1 7465 XNOR2X1 $T=2447280 1723120 0 0 $X=2447278 $Y=1722718
X857 7496 631 3 1 762 XNOR2X1 $T=2461800 1763440 0 0 $X=2461798 $Y=1763038
X858 763 5919 3 1 7578 XNOR2X1 $T=2472360 1622320 1 0 $X=2472358 $Y=1616880
X859 7262 758 3 1 7509 XNOR2X1 $T=2507340 1733200 1 0 $X=2507338 $Y=1727760
X860 776 5936 3 1 7660 XNOR2X1 $T=2512620 1743280 1 0 $X=2512618 $Y=1737840
X861 776 7637 3 1 7781 XNOR2X1 $T=2521860 1702960 0 0 $X=2521858 $Y=1702558
X862 783 6166 3 1 7746 XNOR2X1 $T=2527140 1672720 1 0 $X=2527138 $Y=1667280
X863 7864 633 3 1 788 XNOR2X1 $T=2554860 1662640 0 180 $X=2549580 $Y=1657200
X864 768 767 3 1 7812 XNOR2X1 $T=2556180 1622320 0 0 $X=2556178 $Y=1621918
X865 7703 783 3 1 7897 XNOR2X1 $T=2557500 1672720 1 0 $X=2557498 $Y=1667280
X866 786 7809 3 1 8086 XNOR2X1 $T=2557500 1702960 0 0 $X=2557498 $Y=1702558
X867 7812 791 3 1 7888 XNOR2X1 $T=2559480 1642480 1 0 $X=2559478 $Y=1637040
X868 7825 792 3 1 7898 XNOR2X1 $T=2559480 1702960 1 0 $X=2559478 $Y=1697520
X869 7781 7898 3 1 7963 XNOR2X1 $T=2567400 1702960 1 0 $X=2567398 $Y=1697520
X870 2576 90 3 90 1 2575 2612 109 OAI221XL $T=928620 1713040 0 180 $X=924000 $Y=1707600
X871 227 243 3 240 1 238 3479 3109 OAI221XL $T=1200540 1652560 1 180 $X=1195920 $Y=1652158
X872 227 317 3 314 1 242 3789 321 OAI221XL $T=1286340 1733200 1 0 $X=1286338 $Y=1727760
X873 227 302 3 333 1 238 3875 331 OAI221XL $T=1321980 1733200 0 180 $X=1317360 $Y=1727760
X874 227 340 3 341 1 238 3886 3895 OAI221XL $T=1327920 1733200 0 0 $X=1327918 $Y=1732798
X875 487 601 3 600 1 505 5483 5754 OAI221XL $T=1931820 1632400 0 180 $X=1927200 $Y=1626960
X876 608 505 3 487 1 314 5771 5714 OAI221XL $T=1933800 1753360 0 180 $X=1929180 $Y=1747920
X877 487 323 3 602 1 505 5741 5774 OAI221XL $T=1934460 1733200 1 180 $X=1929840 $Y=1732798
X878 487 333 3 5814 1 533 5756 5802 OAI221XL $T=1938420 1723120 1 180 $X=1933800 $Y=1722718
X879 487 258 3 607 1 505 5505 5842 OAI221XL $T=1950300 1632400 1 180 $X=1945680 $Y=1631998
X880 8043 837 3 837 1 8047 8061 832 OAI221XL $T=2628780 1642480 0 180 $X=2624160 $Y=1637040
X881 37 35 30 1 3 25 ADDHXL $T=689700 1753360 0 180 $X=682440 $Y=1747920
X882 4433 4424 123 1 3 396 ADDHXL $T=1489620 1773520 1 180 $X=1482360 $Y=1773118
X883 420 4583 365 1 3 4433 ADDHXL $T=1537140 1773520 0 180 $X=1529880 $Y=1768080
X884 5022 5020 457 1 3 467 ADDHXL $T=1662540 1773520 0 180 $X=1655280 $Y=1768080
X885 5048 5008 465 1 3 5022 ADDHXL $T=1669800 1723120 1 180 $X=1662540 $Y=1722718
X886 380 5049 456 1 3 5048 ADDHXL $T=1663200 1713040 0 0 $X=1663198 $Y=1712638
X887 7026 6935 718 1 3 6979 ADDHXL $T=2310000 1662640 1 180 $X=2302740 $Y=1662238
X888 7088 7085 718 1 3 725 ADDHXL $T=2337060 1622320 0 180 $X=2329800 $Y=1616880
X889 1 6435 6400 6439 3 NOR2XL $T=2137740 1702960 1 0 $X=2137738 $Y=1697520
X890 1 549 6715 6772 3 NOR2XL $T=2228160 1682800 1 0 $X=2228158 $Y=1677360
X891 1 6844 6858 6799 3 NOR2XL $T=2256540 1743280 1 0 $X=2256538 $Y=1737840
X892 1 544 6784 6889 3 NOR2XL $T=2269740 1672720 1 0 $X=2269738 $Y=1667280
X893 1 7070 726 737 3 NOR2XL $T=2356200 1773520 0 0 $X=2356198 $Y=1773118
X894 1 608 7262 748 3 NOR2XL $T=2399100 1763440 0 0 $X=2399098 $Y=1763038
X895 1 7980 8022 7981 3 NOR2XL $T=2601060 1682800 0 180 $X=2599080 $Y=1677360
X896 6326 6372 6366 3 1 6360 XOR3X2 $T=2125200 1723120 0 180 $X=2113320 $Y=1717680
X897 629 623 668 3 1 665 XOR3X2 $T=2135760 1753360 1 180 $X=2123880 $Y=1752958
X898 621 5936 623 3 1 6622 XOR3X2 $T=2189220 1743280 0 0 $X=2189218 $Y=1742878
X899 6621 6627 6706 3 1 6710 XOR3X2 $T=2206380 1713040 1 0 $X=2206378 $Y=1707600
X900 692 6938 6928 3 1 709 XOR3X2 $T=2292180 1632400 1 180 $X=2280300 $Y=1631998
X901 7511 7411 7479 3 1 759 XOR3X2 $T=2468400 1713040 1 180 $X=2456520 $Y=1712638
X902 5929 633 768 3 1 7556 XOR3X2 $T=2484900 1723120 0 0 $X=2484898 $Y=1722718
X903 7636 773 7635 3 1 7733 XOR3X2 $T=2513940 1632400 0 0 $X=2513938 $Y=1631998
X904 7582 7719 7721 3 1 784 XOR3X2 $T=2517240 1773520 1 0 $X=2517238 $Y=1768080
X905 7697 7800 7804 3 1 7801 XOR3X2 $T=2539680 1682800 0 0 $X=2539678 $Y=1682398
X906 7733 7827 7818 3 1 789 XOR3X2 $T=2542320 1733200 1 0 $X=2542318 $Y=1727760
X907 7801 7815 7836 3 1 793 XOR3X2 $T=2542320 1773520 0 0 $X=2542318 $Y=1773118
X908 7925 7948 7940 3 1 6891 XOR3X2 $T=2592480 1662640 0 180 $X=2580600 $Y=1657200
X909 7777 600 7864 3 1 7948 XOR3X2 $T=2583240 1632400 1 0 $X=2583238 $Y=1626960
X910 6546 6470 1 6549 3 6551 AOI21XL $T=2168760 1652560 1 0 $X=2168758 $Y=1647120
X911 8077 8075 1 8022 3 8055 AOI21XL $T=2616240 1662640 1 180 $X=2613600 $Y=1662238
X912 2576 90 2579 3 2606 1 OAI2BB1X1 $T=915420 1713040 0 0 $X=915418 $Y=1712638
X913 3172 3162 3185 3 3161 1 OAI2BB1X1 $T=1099560 1743280 1 0 $X=1099558 $Y=1737840
X914 418 4582 419 3 4640 1 OAI2BB1X1 $T=1531860 1642480 1 0 $X=1531858 $Y=1637040
X915 448 4736 449 3 4831 1 OAI2BB1X1 $T=1589280 1622320 1 0 $X=1589278 $Y=1616880
X916 6637 6622 608 3 6680 1 OAI2BB1X1 $T=2202420 1763440 0 0 $X=2202418 $Y=1763038
X917 6734 6727 6724 3 693 1 OAI2BB1X1 $T=2222880 1642480 0 180 $X=2219580 $Y=1637040
X918 7023 5814 7050 3 7070 1 OAI2BB1X1 $T=2315280 1763440 1 0 $X=2315278 $Y=1758000
X919 7123 602 7151 3 728 1 OAI2BB1X1 $T=2357520 1743280 1 180 $X=2354220 $Y=1742878
X920 7248 7222 7249 3 741 1 OAI2BB1X1 $T=2391180 1702960 1 180 $X=2387880 $Y=1702558
X921 7260 7301 7257 3 749 1 OAI2BB1X1 $T=2401080 1753360 1 0 $X=2401078 $Y=1747920
X922 7329 7331 7315 3 750 1 OAI2BB1X1 $T=2410980 1753360 0 180 $X=2407680 $Y=1747920
X923 756 633 7348 3 7250 1 OAI2BB1X1 $T=2420220 1642480 1 180 $X=2416920 $Y=1642078
X924 626 621 7466 3 7494 1 OAI2BB1X1 $T=2451240 1662640 0 0 $X=2451238 $Y=1662238
X925 7491 7492 7510 3 777 1 OAI2BB1X1 $T=2469060 1682800 1 0 $X=2469058 $Y=1677360
X926 7511 7479 7411 3 7537 1 OAI2BB1X1 $T=2471700 1713040 1 0 $X=2471698 $Y=1707600
X927 7636 7635 773 3 7641 1 OAI2BB1X1 $T=2503380 1632400 0 0 $X=2503378 $Y=1631998
X928 7556 7587 7638 3 775 1 OAI2BB1X1 $T=2503380 1753360 1 0 $X=2503378 $Y=1747920
X929 768 776 7676 3 7912 1 OAI2BB1X1 $T=2527800 1723120 1 0 $X=2527798 $Y=1717680
X930 7800 7804 7697 3 7837 1 OAI2BB1X1 $T=2542320 1672720 0 0 $X=2542318 $Y=1672318
X931 7801 7836 7816 3 787 1 OAI2BB1X1 $T=2548260 1773520 0 180 $X=2544960 $Y=1768080
X932 7733 7818 7862 3 790 1 OAI2BB1X1 $T=2552880 1723120 0 0 $X=2552878 $Y=1722718
X933 7781 7825 792 3 7887 1 OAI2BB1X1 $T=2560800 1692880 1 0 $X=2560798 $Y=1687440
X934 7701 7703 7900 3 7925 1 OAI2BB1X1 $T=2568720 1662640 1 0 $X=2568718 $Y=1657200
X935 7465 7912 7916 3 796 1 OAI2BB1X1 $T=2575320 1743280 1 0 $X=2575318 $Y=1737840
X936 7931 797 7644 3 7941 1 OAI2BB1X1 $T=2585220 1743280 1 180 $X=2581920 $Y=1742878
X937 7864 7777 600 3 7952 1 OAI2BB1X1 $T=2584560 1642480 1 0 $X=2584558 $Y=1637040
X938 7509 803 7990 3 8059 1 OAI2BB1X1 $T=2599080 1723120 0 0 $X=2599078 $Y=1722718
X939 8094 8022 8074 3 8080 1 OAI2BB1X1 $T=2620200 1652560 0 180 $X=2616900 $Y=1647120
X940 8086 8059 8093 3 8095 1 OAI2BB1X1 $T=2619540 1702960 0 0 $X=2619538 $Y=1702558
X941 1896 3 1915 1 1962 NAND2BXL $T=713460 1662640 0 0 $X=713458 $Y=1662238
X942 2080 3 2005 1 2104 NAND2BXL $T=762960 1692880 1 0 $X=762958 $Y=1687440
X943 2118 3 2112 1 2106 NAND2BXL $T=774840 1672720 1 180 $X=772200 $Y=1672318
X944 89 3 34 1 2540 NAND2BXL $T=906840 1733200 0 180 $X=904200 $Y=1727760
X945 2493 3 2516 1 2590 NAND2BXL $T=914760 1692880 1 0 $X=914758 $Y=1687440
X946 3210 3 3152 1 3122 NAND2BXL $T=1096260 1632400 1 180 $X=1093620 $Y=1631998
X947 3963 3 3954 1 3898 NAND2BXL $T=1346400 1672720 1 180 $X=1343760 $Y=1672318
X948 3990 3 4010 1 3948 NAND2BXL $T=1362240 1662640 0 180 $X=1359600 $Y=1657200
X949 7550 3 631 1 7809 NAND2BXL $T=2539020 1702960 0 0 $X=2539018 $Y=1702558
X950 73 69 75 2302 1 3 77 AOI2BB2X1 $T=827640 1773520 0 0 $X=827638 $Y=1773118
X951 3297 211 213 215 1 3 3418 AOI2BB2X1 $T=1171500 1632400 0 0 $X=1171498 $Y=1631998
X952 218 219 222 226 1 3 224 AOI2BB2X1 $T=1184700 1632400 0 0 $X=1184698 $Y=1631998
X953 3516 219 245 226 1 3 3488 AOI2BB2X1 $T=1203180 1723120 1 180 $X=1198560 $Y=1722718
X954 304 219 320 283 1 3 3789 AOI2BB2X1 $T=1286340 1733200 0 0 $X=1286338 $Y=1732798
X955 281 3664 329 226 1 3 3875 AOI2BB2X1 $T=1307460 1733200 1 0 $X=1307458 $Y=1727760
X956 492 5276 220 493 1 3 5302 AOI2BB2X1 $T=1746360 1713040 1 0 $X=1746358 $Y=1707600
X957 494 5276 234 493 1 3 5259 AOI2BB2X1 $T=1751640 1692880 1 180 $X=1747020 $Y=1692478
X958 496 5276 213 493 1 3 5308 AOI2BB2X1 $T=1758240 1692880 1 180 $X=1753620 $Y=1692478
X959 513 510 236 493 1 3 5371 AOI2BB2X1 $T=1784640 1642480 0 180 $X=1780020 $Y=1637040
X960 517 510 493 230 1 3 5406 AOI2BB2X1 $T=1795860 1642480 0 180 $X=1791240 $Y=1637040
X961 531 5276 493 245 1 3 5509 AOI2BB2X1 $T=1813680 1713040 1 0 $X=1813678 $Y=1707600
X962 5500 510 493 222 1 3 5483 AOI2BB2X1 $T=1820940 1642480 0 180 $X=1816320 $Y=1637040
X963 542 5276 493 300 1 3 5488 AOI2BB2X1 $T=1822260 1733200 0 180 $X=1817640 $Y=1727760
X964 546 510 221 493 1 3 5505 AOI2BB2X1 $T=1826880 1632400 1 180 $X=1822260 $Y=1631998
X965 572 5276 493 287 1 3 5551 AOI2BB2X1 $T=1849320 1733200 1 180 $X=1844700 $Y=1732798
X966 587 5276 336 493 1 3 5766 AOI2BB2X1 $T=1896180 1743280 0 0 $X=1896178 $Y=1742878
X967 592 5276 324 493 1 3 5741 AOI2BB2X1 $T=1907400 1733200 0 0 $X=1907398 $Y=1732798
X968 591 5276 320 493 1 3 5771 AOI2BB2X1 $T=1907400 1753360 1 0 $X=1907398 $Y=1747920
X969 593 5276 493 329 1 3 5756 AOI2BB2X1 $T=1908720 1723120 0 0 $X=1908718 $Y=1722718
X970 2274 3 2273 1 2272 2181 NAND3X1 $T=821700 1652560 0 180 $X=819060 $Y=1647120
X971 2393 3 2392 1 2391 2336 NAND3X1 $T=858660 1662640 0 180 $X=856020 $Y=1657200
X972 3418 3 3406 1 3481 3113 NAND3X1 $T=1174800 1642480 0 180 $X=1172160 $Y=1637040
X973 3436 3 3437 1 3438 2748 NAND3X1 $T=1184040 1632400 1 0 $X=1184038 $Y=1626960
X974 3461 3 3468 1 3471 3425 NAND3X1 $T=1194600 1682800 0 0 $X=1194598 $Y=1682398
X975 365 3 130 1 123 4437 NAND3X1 $T=1503480 1733200 0 180 $X=1500840 $Y=1727760
X976 4528 3 130 1 123 4432 NAND3X1 $T=1513380 1733200 1 180 $X=1510740 $Y=1732798
X977 4598 3 4599 1 4601 4337 NAND3X1 $T=1539120 1692880 1 0 $X=1539118 $Y=1687440
X978 4927 3 457 1 464 4872 NAND3X1 $T=1639440 1763440 0 180 $X=1636800 $Y=1758000
X979 4949 3 4971 1 4911 4832 NAND3X1 $T=1642080 1743280 0 180 $X=1639440 $Y=1737840
X980 5009 3 5010 1 4979 5018 NAND3X1 $T=1653300 1702960 1 0 $X=1653298 $Y=1697520
X981 380 3 5038 1 4975 5050 NAND3X1 $T=1662540 1692880 0 0 $X=1662538 $Y=1692478
X982 5309 3 5311 1 5308 5334 NAND3X1 $T=1755600 1682800 0 0 $X=1755598 $Y=1682398
X983 5758 3 5766 1 5768 596 NAND3X1 $T=1919280 1753360 0 0 $X=1919278 $Y=1752958
X984 8020 3 8075 1 8094 837 NAND3X1 $T=2628120 1642480 0 0 $X=2628118 $Y=1642078
X985 5919 633 614 6608 3 1 6564 CMPR32X1 $T=2201760 1692880 0 180 $X=2187900 $Y=1687440
X986 6937 7043 6971 3 7017 1 AOI2BB1X2 $T=2306040 1692880 1 180 $X=2301420 $Y=1692478
X987 404 423 3 1 4612 OR2X1 $T=1541100 1622320 1 0 $X=1541098 $Y=1616880
X988 53 1 45 3 CLKINVX3 $T=728640 1632400 0 180 $X=726660 $Y=1626960
X989 1999 1 2027 3 CLKINVX3 $T=742500 1723120 0 0 $X=742498 $Y=1722718
X990 2109 1 2094 3 CLKINVX3 $T=773520 1662640 1 0 $X=773518 $Y=1657200
X991 86 1 2382 3 CLKINVX3 $T=867900 1692880 1 0 $X=867898 $Y=1687440
X992 94 1 2422 3 CLKINVX3 $T=889020 1733200 0 180 $X=887040 $Y=1727760
X993 2966 1 2900 3 CLKINVX3 $T=1032900 1743280 1 0 $X=1032898 $Y=1737840
X994 89 1 171 3 CLKINVX3 $T=1075800 1753360 1 0 $X=1075798 $Y=1747920
X995 245 1 249 3 CLKINVX3 $T=1209120 1733200 0 0 $X=1209118 $Y=1732798
X996 3719 1 301 3 CLKINVX3 $T=1261260 1692880 0 0 $X=1261258 $Y=1692478
X997 325 1 3784 3 CLKINVX3 $T=1301520 1652560 0 0 $X=1301518 $Y=1652158
X998 3842 1 3664 3 CLKINVX3 $T=1312740 1702960 0 0 $X=1312738 $Y=1702558
X999 4512 1 4436 3 CLKINVX3 $T=1512720 1733200 1 0 $X=1512718 $Y=1727760
X1000 428 1 451 3 CLKINVX3 $T=1593240 1763440 0 0 $X=1593238 $Y=1763038
X1001 4833 1 4835 3 CLKINVX3 $T=1602480 1672720 1 0 $X=1602478 $Y=1667280
X1002 473 1 240 3 CLKINVX3 $T=1679040 1682800 0 0 $X=1679038 $Y=1682398
X1003 5267 1 492 3 CLKINVX3 $T=1740420 1713040 0 180 $X=1738440 $Y=1707600
X1004 485 1 494 3 CLKINVX3 $T=1750980 1773520 0 0 $X=1750978 $Y=1773118
X1005 492 1 501 3 CLKINVX3 $T=1778700 1702960 1 0 $X=1778698 $Y=1697520
X1006 518 1 531 3 CLKINVX3 $T=1815000 1692880 0 0 $X=1814998 $Y=1692478
X1007 575 1 563 3 CLKINVX3 $T=1853280 1713040 0 180 $X=1851300 $Y=1707600
X1008 5757 1 593 3 CLKINVX3 $T=1913340 1662640 0 180 $X=1911360 $Y=1657200
X1009 5978 1 607 3 CLKINVX3 $T=2055240 1632400 0 180 $X=2053260 $Y=1626960
X1010 629 1 5814 3 CLKINVX3 $T=2112660 1763440 1 0 $X=2112658 $Y=1758000
X1011 633 1 5920 3 CLKINVX3 $T=2173380 1733200 0 0 $X=2173378 $Y=1732798
X1012 5814 1 6342 3 CLKINVX3 $T=2196480 1753360 0 0 $X=2196478 $Y=1752958
X1013 544 1 557 3 CLKINVX3 $T=2233440 1743280 1 180 $X=2231460 $Y=1742878
X1014 536 1 561 3 CLKINVX3 $T=2273040 1692880 1 0 $X=2273038 $Y=1687440
X1015 605 1 718 3 CLKINVX3 $T=2363460 1702960 0 180 $X=2361480 $Y=1697520
X1016 5919 1 754 3 CLKINVX3 $T=2416260 1632400 1 0 $X=2416258 $Y=1626960
X1017 6166 1 727 3 CLKINVX3 $T=2420220 1662640 1 0 $X=2420218 $Y=1657200
X1018 626 1 613 3 CLKINVX3 $T=2445300 1622320 1 0 $X=2445298 $Y=1616880
X1019 5936 1 756 3 CLKINVX3 $T=2463780 1642480 0 0 $X=2463778 $Y=1642078
X1020 5929 1 758 3 CLKINVX3 $T=2494800 1682800 0 0 $X=2494798 $Y=1682398
X1021 443 426 1 3 356 AND2X1 $T=1584000 1662640 1 0 $X=1583998 $Y=1657200
X1022 6250 6255 1 3 6248 AND2X1 $T=2088900 1642480 1 180 $X=2086260 $Y=1642078
X1023 6932 6937 1 3 6947 AND2X1 $T=2284920 1713040 1 0 $X=2284918 $Y=1707600
X1024 34 193 1 194 195 3289 3 AOI22X1 $T=1134540 1763440 1 0 $X=1134538 $Y=1758000
X1025 199 194 1 196 94 3296 3 AOI22X1 $T=1141140 1723120 0 0 $X=1141138 $Y=1722718
X1026 4567 410 1 415 421 4556 3 AOI22X1 $T=1535820 1753360 1 0 $X=1535818 $Y=1747920
X1027 4662 428 1 427 425 4549 3 AOI22X1 $T=1554300 1763440 1 180 $X=1551000 $Y=1763038
X1028 543 5393 1 506 500 5529 3 AOI22X1 $T=1830840 1682800 0 0 $X=1830838 $Y=1682398
X1029 8056 8096 1 8096 805 8083 3 AOI22X1 $T=2626140 1662640 0 180 $X=2622840 $Y=1657200
X1030 482 476 476 4971 3 1 5155 OAI2BB2X1 $T=1705440 1753360 1 180 $X=1700820 $Y=1752958
X1031 480 476 476 4911 3 1 5156 OAI2BB2X1 $T=1706760 1743280 0 180 $X=1702140 $Y=1737840
X1032 481 476 476 5070 3 1 5181 OAI2BB2X1 $T=1710060 1692880 1 0 $X=1710058 $Y=1687440
X1033 6262 605 6290 649 3 1 6326 OAI2BB2X1 $T=2095500 1753360 1 0 $X=2095498 $Y=1747920
X1034 730 728 733 7112 3 1 735 OAI2BB2X1 $T=2348940 1773520 1 0 $X=2348938 $Y=1768080
X1035 551 561 3 1 6627 XNOR2XL $T=2201100 1702960 1 0 $X=2201098 $Y=1697520
X1036 557 576 3 1 6795 XNOR2XL $T=2228160 1753360 0 0 $X=2228158 $Y=1752958
X1037 578 535 3 1 6855 XNOR2XL $T=2240700 1773520 1 0 $X=2240698 $Y=1768080
X1038 544 6859 3 1 705 XNOR2XL $T=2256540 1632400 1 0 $X=2256538 $Y=1626960
X1039 613 772 3 1 7701 XNOR2XL $T=2545620 1632400 1 0 $X=2545618 $Y=1626960
X1040 2154 99 2476 1 3 OR2X4 $T=886380 1632400 1 0 $X=886378 $Y=1626960
X1041 3784 3770 207 1 3 OR2X4 $T=1285680 1642480 1 180 $X=1281720 $Y=1642078
X1042 3784 316 212 1 3 OR2X4 $T=1288320 1652560 1 180 $X=1284360 $Y=1652158
X1043 3784 316 202 1 3 OR2X4 $T=1296900 1652560 1 0 $X=1296898 $Y=1647120
X1044 3842 3868 242 1 3 OR2X4 $T=1314060 1642480 1 0 $X=1314058 $Y=1637040
X1045 2620 353 4077 1 3 OR2X4 $T=1380720 1622320 0 0 $X=1380718 $Y=1621918
X1046 4799 4927 4931 1 3 OR2X4 $T=1630860 1723120 0 0 $X=1630858 $Y=1722718
X1047 5303 3868 5275 1 3 OR2X4 $T=1753620 1642480 0 180 $X=1749660 $Y=1637040
X1048 5303 3770 505 1 3 OR2X4 $T=1772760 1632400 0 0 $X=1772758 $Y=1631998
X1049 5757 5767 599 1 3 OR2X4 $T=1927200 1652560 0 0 $X=1927198 $Y=1652158
X1050 619 5958 617 1 3 OR2X4 $T=1991880 1702960 0 180 $X=1987920 $Y=1697520
X1051 2027 49 1963 3 1 2142 OAI2BB1X4 $T=755700 1723120 1 0 $X=755698 $Y=1717680
X1052 392 123 4380 3 1 4387 OAI2BB1X4 $T=1469820 1763440 1 0 $X=1469818 $Y=1758000
X1053 394 4396 4365 3 1 4350 OAI2BB1X4 $T=1477740 1733200 0 180 $X=1471140 $Y=1727760
X1054 4590 418 419 3 1 401 OAI2BB1X4 $T=1536480 1652560 0 180 $X=1529880 $Y=1647120
X1055 3605 285 3 1 INVX8 $T=1239480 1773520 1 0 $X=1239478 $Y=1768080
X1056 3844 227 3 1 INVX8 $T=1306800 1632400 1 180 $X=1302840 $Y=1631998
X1057 4471 403 3 1 INVX8 $T=1498200 1682800 1 0 $X=1498198 $Y=1677360
X1058 4463 417 3 1 INVX8 $T=1508760 1622320 1 0 $X=1508758 $Y=1616880
X1059 352 316 3 1 INVX8 $T=1514040 1652560 0 0 $X=1514038 $Y=1652158
X1060 4686 4512 3 1 INVX8 $T=1564200 1632400 1 0 $X=1564198 $Y=1626960
X1061 4868 428 3 1 INVX8 $T=1618320 1652560 0 0 $X=1618318 $Y=1652158
X1062 654 608 3 1 INVX8 $T=2092200 1773520 1 0 $X=2092198 $Y=1768080
X1063 6353 5936 3 1 INVX8 $T=2285580 1723120 1 0 $X=2285578 $Y=1717680
X1064 61 2082 1999 3 1 NAND2BX2 $T=764280 1763440 0 180 $X=760320 $Y=1758000
X1065 2587 4025 4065 3 1 NAND2BX2 $T=1366860 1642480 0 0 $X=1366858 $Y=1642078
X1066 49 1989 1982 1961 1 3 OAI2BB1X2 $T=739200 1713040 0 180 $X=734580 $Y=1707600
X1067 2809 2808 2804 129 1 3 OAI2BB1X2 $T=992640 1632400 1 180 $X=988020 $Y=1631998
X1068 3132 3161 3165 3167 1 3 OAI2BB1X2 $T=1095600 1702960 0 0 $X=1095598 $Y=1702558
X1069 393 4365 4356 4323 1 3 OAI2BB1X2 $T=1467180 1753360 0 180 $X=1462560 $Y=1747920
X1070 4463 404 402 4476 1 3 OAI2BB1X2 $T=1502820 1622320 0 180 $X=1498200 $Y=1616880
X1071 506 512 5390 515 1 3 OAI2BB1X2 $T=1785300 1763440 0 0 $X=1785298 $Y=1763038
X1072 812 8073 813 3 1 8045 AND3X1 $T=2614920 1632400 0 180 $X=2611620 $Y=1626960
X1073 8075 8073 8094 3 1 8096 AND3X1 $T=2629440 1652560 1 180 $X=2626140 $Y=1652158
X1074 4927 4971 457 3 1 4985 AND3X2 $T=1646700 1753360 1 0 $X=1646698 $Y=1747920
X1075 456 380 465 3 1 4927 AND3X2 $T=1656600 1723120 1 180 $X=1653300 $Y=1722718
X1076 4641 4658 4598 3 1 NOR2BX2 $T=1550340 1642480 0 0 $X=1550338 $Y=1642078
X1077 7493 7495 761 3 1 NOR2BX2 $T=2461140 1733200 0 0 $X=2461138 $Y=1732798
X1078 30 29 3 1 24 XOR2XL $T=673860 1662640 1 180 $X=668580 $Y=1662238
X1079 632 602 3 1 7496 XOR2XL $T=2434080 1763440 1 0 $X=2434078 $Y=1758000
X1080 1 3462 2780 3454 3450 3 NAND3X2 $T=1187340 1723120 0 0 $X=1187338 $Y=1722718
X1081 1 377 4171 4264 4272 3 NAND3X2 $T=1442760 1773520 1 180 $X=1438140 $Y=1773118
X1082 1 4322 4243 4321 385 3 NAND3X2 $T=1448700 1773520 1 0 $X=1448698 $Y=1768080
X1083 1 4340 4255 4325 388 3 NAND3X2 $T=1450680 1743280 0 0 $X=1450678 $Y=1742878
X1084 1 4351 4338 4350 4272 3 NAND3X2 $T=1459260 1733200 1 0 $X=1459258 $Y=1727760
X1085 1 4349 4326 4370 4272 3 NAND3X2 $T=1459260 1743280 0 0 $X=1459258 $Y=1742878
X1086 1 4549 4372 4540 4556 3 NAND3X2 $T=1523280 1753360 0 180 $X=1518660 $Y=1747920
X1087 1 4944 462 4929 4871 3 NAND3X2 $T=1632840 1753360 0 0 $X=1632838 $Y=1752958
X1088 118 117 125 2728 112 1 3 2670 SDFFRHQXL $T=972840 1723120 0 180 $X=956340 $Y=1717680
X1089 118 117 126 2748 112 1 3 2715 SDFFRHQXL $T=974160 1632400 0 180 $X=957660 $Y=1626960
X1090 118 117 119 2731 112 1 3 2662 SDFFRHQXL $T=974160 1652560 1 180 $X=957660 $Y=1652158
X1091 118 117 114 2756 112 1 3 2703 SDFFRHQXL $T=975480 1702960 0 180 $X=958980 $Y=1697520
X1092 118 117 110 2732 112 1 3 2716 SDFFRHQXL $T=959640 1672720 0 0 $X=959638 $Y=1672318
X1093 118 117 27 3000 112 1 3 2935 SDFFRHQXL $T=1055340 1632400 0 180 $X=1038840 $Y=1626960
X1094 118 117 89 159 112 1 3 2989 SDFFRHQXL $T=1055340 1642480 0 180 $X=1038840 $Y=1637040
X1095 118 117 29 3134 112 1 3 173 SDFFRHQXL $T=1094940 1622320 1 180 $X=1078440 $Y=1621918
X1096 118 117 276 3626 291 1 3 3639 SDFFRHQXL $T=1230240 1652560 0 0 $X=1230238 $Y=1652158
X1097 118 117 293 3728 169 1 3 3733 SDFFRHQXL $T=1262580 1672720 0 0 $X=1262578 $Y=1672318
X1098 364 117 157 4171 169 1 3 358 SDFFRHQXL $T=1409100 1773520 0 180 $X=1392600 $Y=1768080
X1099 364 117 130 4243 169 1 3 4195 SDFFRHQXL $T=1439460 1773520 0 180 $X=1422960 $Y=1768080
X1100 364 117 365 4255 169 1 3 4180 SDFFRHQXL $T=1442100 1743280 0 180 $X=1425600 $Y=1737840
X1101 364 117 380 4260 169 1 3 4206 SDFFRHQXL $T=1444080 1733200 0 180 $X=1427580 $Y=1727760
X1102 364 117 386 4326 169 1 3 4366 SDFFRHQXL $T=1450680 1723120 0 0 $X=1450678 $Y=1722718
X1103 364 117 122 4335 169 1 3 4348 SDFFRHQXL $T=1453980 1672720 1 0 $X=1453978 $Y=1667280
X1104 364 117 387 4337 169 1 3 4379 SDFFRHQXL $T=1454640 1682800 1 0 $X=1454638 $Y=1677360
X1105 364 117 123 4338 169 1 3 4364 SDFFRHQXL $T=1454640 1702960 1 0 $X=1454638 $Y=1697520
X1106 364 478 480 5155 483 1 3 5179 SDFFRHQXL $T=1696200 1753360 1 0 $X=1696198 $Y=1747920
X1107 364 479 481 5011 483 1 3 456 SDFFRHQXL $T=1698840 1652560 0 0 $X=1698838 $Y=1652158
X1108 364 479 456 5072 483 1 3 5167 SDFFRHQXL $T=1698840 1682800 1 0 $X=1698838 $Y=1677360
X1109 364 479 465 5156 483 1 3 5189 SDFFRHQXL $T=1698840 1713040 0 0 $X=1698838 $Y=1712638
X1110 364 479 488 5181 483 1 3 5165 SDFFRHQXL $T=1735140 1632400 1 180 $X=1718640 $Y=1631998
X1111 364 478 490 5235 491 1 3 5267 SDFFRHQXL $T=1730520 1713040 0 0 $X=1730518 $Y=1712638
X1112 364 478 500 5335 491 1 3 495 SDFFRHQXL $T=1769460 1773520 0 180 $X=1752960 $Y=1768080
X1113 364 479 504 5359 483 1 3 5386 SDFFRHQXL $T=1768800 1672720 0 0 $X=1768798 $Y=1672318
X1114 364 478 507 5373 491 1 3 525 SDFFRHQXL $T=1776060 1753360 1 0 $X=1776058 $Y=1747920
X1115 364 478 540 5506 491 1 3 500 SDFFRHQXL $T=1827540 1763440 1 180 $X=1811040 $Y=1763038
X1116 364 478 556 5550 491 1 3 552 SDFFRHQXL $T=1876380 1743280 0 180 $X=1859880 $Y=1737840
X1117 364 478 580 5560 491 1 3 5635 SDFFRHQXL $T=1860540 1702960 1 0 $X=1860538 $Y=1697520
X1118 364 478 552 5616 491 1 3 5636 SDFFRHQXL $T=1860540 1733200 1 0 $X=1860538 $Y=1727760
X1119 364 478 582 583 491 1 3 556 SDFFRHQXL $T=1862520 1773520 1 0 $X=1862518 $Y=1768080
X1120 364 478 536 570 491 1 3 5715 SDFFRHQXL $T=1886280 1632400 1 0 $X=1886278 $Y=1626960
X1121 364 478 574 5754 491 1 3 5726 SDFFRHQXL $T=1921260 1632400 1 180 $X=1904760 $Y=1631998
X1122 364 478 594 5842 491 1 3 5876 SDFFRHQXL $T=1943040 1642480 0 0 $X=1943038 $Y=1642078
X1123 364 478 5973 5970 491 1 3 6015 SDFFRHQXL $T=1989240 1672720 1 0 $X=1989238 $Y=1667280
X1124 364 478 5978 5928 491 1 3 6020 SDFFRHQXL $T=1991880 1622320 0 0 $X=1991878 $Y=1621918
X1125 364 588 621 5927 491 1 3 6046 SDFFRHQXL $T=1993200 1733200 0 0 $X=1993198 $Y=1732798
X1126 364 588 623 5926 491 1 3 6059 SDFFRHQXL $T=1993860 1723120 0 0 $X=1993858 $Y=1722718
X1127 364 588 620 5980 491 1 3 6028 SDFFRHQXL $T=1994520 1763440 1 0 $X=1994518 $Y=1758000
X1128 364 478 6048 5957 491 1 3 6096 SDFFRHQXL $T=2014320 1672720 1 0 $X=2014318 $Y=1667280
X1129 364 478 631 5935 491 1 3 6048 SDFFRHQXL $T=2014320 1672720 0 0 $X=2014318 $Y=1672318
X1130 364 478 632 6044 491 1 3 5978 SDFFRHQXL $T=2016960 1632400 0 0 $X=2016958 $Y=1631998
X1131 364 478 6055 5918 491 1 3 6128 SDFFRHQXL $T=2016960 1642480 0 0 $X=2016958 $Y=1642078
X1132 364 478 634 5930 491 1 3 636 SDFFRHQXL $T=2018280 1622320 1 0 $X=2018278 $Y=1616880
X1133 97 1 96 3 BUFX3 $T=881100 1743280 0 180 $X=878460 $Y=1737840
X1134 2662 1 110 3 BUFX3 $T=944460 1662640 0 180 $X=941820 $Y=1657200
X1135 2670 1 111 3 BUFX3 $T=947100 1723120 0 180 $X=944460 $Y=1717680
X1136 2716 1 114 3 BUFX3 $T=952380 1672720 1 180 $X=949740 $Y=1672318
X1137 2703 1 115 3 BUFX3 $T=952380 1702960 1 180 $X=949740 $Y=1702558
X1138 2935 1 144 3 BUFX3 $T=1021680 1622320 1 180 $X=1019040 $Y=1621918
X1139 163 1 165 3 BUFX3 $T=1063260 1713040 1 0 $X=1063258 $Y=1707600
X1140 208 1 94 3 BUFX3 $T=1137180 1672720 1 180 $X=1134540 $Y=1672318
X1141 225 1 210 3 BUFX3 $T=1186680 1773520 1 180 $X=1184040 $Y=1773118
X1142 155 1 286 3 BUFX3 $T=1240140 1743280 1 0 $X=1240138 $Y=1737840
X1143 169 1 291 3 BUFX3 $T=1255980 1632400 0 180 $X=1253340 $Y=1626960
X1144 332 1 211 3 BUFX3 $T=1304820 1622320 1 180 $X=1302180 $Y=1621918
X1145 4180 1 130 3 BUFX3 $T=1405800 1743280 0 180 $X=1403160 $Y=1737840
X1146 4206 1 365 3 BUFX3 $T=1411080 1733200 0 180 $X=1408440 $Y=1727760
X1147 4195 1 157 3 BUFX3 $T=1415040 1763440 1 180 $X=1412400 $Y=1763038
X1148 376 1 124 3 BUFX3 $T=1432860 1672720 1 180 $X=1430220 $Y=1672318
X1149 4364 1 122 3 BUFX3 $T=1459920 1692880 0 180 $X=1457280 $Y=1687440
X1150 4348 1 387 3 BUFX3 $T=1460580 1662640 1 180 $X=1457940 $Y=1662238
X1151 4366 1 123 3 BUFX3 $T=1466520 1713040 1 180 $X=1463880 $Y=1712638
X1152 4379 1 380 3 BUFX3 $T=1467840 1692880 0 180 $X=1465200 $Y=1687440
X1153 424 1 4514 3 BUFX3 $T=1605120 1662640 1 0 $X=1605118 $Y=1657200
X1154 474 1 476 3 BUFX3 $T=1680360 1692880 1 0 $X=1680358 $Y=1687440
X1155 5167 1 465 3 BUFX3 $T=1702800 1692880 0 180 $X=1700160 $Y=1687440
X1156 5179 1 482 3 BUFX3 $T=1704120 1763440 1 180 $X=1701480 $Y=1763038
X1157 5165 1 481 3 BUFX3 $T=1709400 1632400 1 180 $X=1706760 $Y=1631998
X1158 478 1 479 3 BUFX3 $T=1718640 1713040 0 180 $X=1716000 $Y=1707600
X1159 5189 1 480 3 BUFX3 $T=1717320 1733200 1 0 $X=1717318 $Y=1727760
X1160 497 1 5276 3 BUFX3 $T=1760880 1642480 1 0 $X=1760878 $Y=1637040
X1161 5386 1 489 3 BUFX3 $T=1783320 1662640 1 180 $X=1780680 $Y=1662238
X1162 497 1 510 3 BUFX3 $T=1790580 1622320 1 0 $X=1790578 $Y=1616880
X1163 5635 1 551 3 BUFX3 $T=1861860 1692880 1 180 $X=1859220 $Y=1692478
X1164 5636 1 580 3 BUFX3 $T=1870440 1723120 0 180 $X=1867800 $Y=1717680
X1165 5726 1 594 3 BUFX3 $T=1906740 1642480 1 0 $X=1906738 $Y=1637040
X1166 5757 1 597 3 BUFX3 $T=1922580 1692880 1 0 $X=1922578 $Y=1687440
X1167 5876 1 543 3 BUFX3 $T=1952940 1642480 0 180 $X=1950300 $Y=1637040
X1168 6020 1 626 3 BUFX3 $T=2003760 1632400 0 180 $X=2001120 $Y=1626960
X1169 6128 1 632 3 BUFX3 $T=2051940 1642480 0 0 $X=2051938 $Y=1642078
X1170 6166 1 5933 3 BUFX3 $T=2057880 1692880 0 0 $X=2057878 $Y=1692478
X1171 5975 1 6353 3 BUFX3 $T=2107380 1713040 1 0 $X=2107378 $Y=1707600
X1172 654 1 6507 3 BUFX3 $T=2152260 1773520 1 0 $X=2152258 $Y=1768080
X1173 4508 4525 1 3 CLKINVX4 $T=1508760 1773520 0 0 $X=1508758 $Y=1773118
X1174 4522 4438 1 3 CLKINVX4 $T=1514040 1743280 1 180 $X=1511400 $Y=1742878
X1175 4728 4562 1 3 CLKINVX4 $T=1576740 1733200 0 180 $X=1574100 $Y=1727760
X1176 4581 4782 1 3 CLKINVX4 $T=1584000 1672720 0 0 $X=1583998 $Y=1672318
X1177 4947 4944 1 3 CLKINVX4 $T=1639440 1753360 0 180 $X=1636800 $Y=1747920
X1178 5202 491 1 3 CLKINVX4 $T=1740420 1763440 0 0 $X=1740418 $Y=1763038
X1179 5467 517 1 3 CLKINVX4 $T=1815000 1672720 1 0 $X=1814998 $Y=1667280
X1180 6048 5929 1 3 CLKINVX4 $T=2034780 1662640 0 0 $X=2034778 $Y=1662238
X1181 28 193 1 196 90 205 194 206 3 AOI222X2 $T=1139820 1622320 1 0 $X=1139818 $Y=1616880
X1182 428 4586 1 421 4512 415 365 4609 3 AOI222X2 $T=1554960 1743280 1 180 $X=1545720 $Y=1742878
X1183 5393 574 1 506 525 5596 575 5383 3 AOI222X2 $T=1849320 1682800 0 0 $X=1849318 $Y=1682398
X1184 604 605 3 341 606 1 603 OAI22X1 $T=1943040 1763440 0 0 $X=1943038 $Y=1763038
X1185 602 604 3 606 323 1 6016 OAI22X1 $T=1970760 1763440 1 180 $X=1966800 $Y=1763038
X1186 5900 604 3 606 251 1 5970 OAI22X1 $T=1973400 1662640 1 180 $X=1969440 $Y=1662238
X1187 613 604 3 606 612 1 5928 OAI22X1 $T=1976040 1622320 0 180 $X=1972080 $Y=1616880
X1188 614 604 3 606 309 1 5980 OAI22X1 $T=1977360 1753360 0 180 $X=1973400 $Y=1747920
X1189 610 604 3 606 615 1 5918 OAI22X1 $T=1980000 1642480 1 180 $X=1976040 $Y=1642078
X1190 607 604 3 606 258 1 6044 OAI22X1 $T=1981320 1632400 1 180 $X=1977360 $Y=1631998
X1191 5919 604 3 606 260 1 5957 OAI22X1 $T=1981320 1672720 0 180 $X=1977360 $Y=1667280
X1192 5929 604 3 606 240 1 5935 OAI22X1 $T=1981320 1672720 1 180 $X=1977360 $Y=1672318
X1193 5933 604 3 606 244 1 5974 OAI22X1 $T=1981320 1702960 1 180 $X=1977360 $Y=1702558
X1194 5936 604 3 606 272 1 6056 OAI22X1 $T=1981320 1713040 1 180 $X=1977360 $Y=1712638
X1195 5920 604 3 606 262 1 5926 OAI22X1 $T=1981320 1723120 1 180 $X=1977360 $Y=1722718
X1196 5921 604 3 606 289 1 5927 OAI22X1 $T=1981320 1733200 1 180 $X=1977360 $Y=1732798
X1197 5814 604 3 606 333 1 616 OAI22X1 $T=1981320 1763440 0 180 $X=1977360 $Y=1758000
X1198 600 604 3 606 601 1 5930 OAI22X1 $T=1983960 1622320 0 180 $X=1980000 $Y=1616880
X1199 730 728 3 726 7070 1 738 OAI22X1 $T=2365440 1773520 1 180 $X=2361480 $Y=1773118
X1200 89 1 34 2543 3 NOR2BXL $T=888360 1702960 0 0 $X=888358 $Y=1702558
X1201 552 1 551 5566 3 NOR2BXL $T=1840740 1713040 0 0 $X=1840738 $Y=1712638
X1202 500 1 576 5531 3 NOR2BXL $T=1855260 1773520 0 0 $X=1855258 $Y=1773118
X1203 556 1 548 5534 3 5531 547 AOI211X1 $T=1836780 1773520 1 180 $X=1833480 $Y=1773118
X1204 3613 273 274 3 210 268 1 275 OAI32X1 $T=1230900 1753360 0 0 $X=1230898 $Y=1752958
X1205 5566 525 563 3 552 560 1 5561 OAI32X1 $T=1848000 1723120 1 180 $X=1843380 $Y=1722718
X1206 5531 556 548 3 500 564 1 5556 OAI32X1 $T=1849320 1773520 1 180 $X=1844700 $Y=1773118
X1207 2576 2575 3 1 2608 2612 AOI2BB1X1 $T=923340 1723120 1 0 $X=923338 $Y=1717680
X1208 262 487 3 1 5841 5516 AOI2BB1X1 $T=1948320 1713040 1 180 $X=1945020 $Y=1712638
X1209 309 487 3 1 5845 5609 AOI2BB1X1 $T=1947660 1723120 0 0 $X=1947658 $Y=1722718
X1210 289 487 3 1 5847 5729 AOI2BB1X1 $T=1948980 1733200 0 0 $X=1948978 $Y=1732798
X1211 767 766 3 1 7579 7636 AOI2BB1X1 $T=2491500 1632400 0 0 $X=2491498 $Y=1631998
X1212 7864 7777 3 1 600 7923 AOI2BB1X1 $T=2576640 1632400 0 0 $X=2576638 $Y=1631998
X1213 520 509 1 506 495 489 5332 508 3 AOI222X1 $T=1783980 1773520 1 180 $X=1778700 $Y=1773118
X1214 559 5393 1 506 552 551 5541 509 3 AOI222X1 $T=1844700 1682800 1 180 $X=1839420 $Y=1682398
X1215 778 811 1 812 8058 8056 810 8045 3 AOI222X1 $T=2609640 1622320 1 0 $X=2609638 $Y=1616880
X1216 7777 7864 3 7888 1 7952 8020 OAI211X1 $T=2583900 1642480 0 0 $X=2583898 $Y=1642078
X1217 8055 8081 3 8083 1 8074 8023 OAI211X1 $T=2615580 1662640 1 0 $X=2615578 $Y=1657200
X1218 6262 605 649 3 1 6214 XNOR3X2 $T=2089560 1753360 1 180 $X=2077680 $Y=1752958
X1219 7023 7013 6976 3 1 715 XNOR3X2 $T=2306700 1733200 1 180 $X=2294820 $Y=1732798
X1220 7123 7191 7185 3 1 726 XNOR3X2 $T=2364780 1743280 0 0 $X=2364778 $Y=1742878
X1221 7260 6166 7301 3 1 7331 XNOR3X2 $T=2402400 1743280 1 0 $X=2402398 $Y=1737840
X1222 7556 7444 7587 3 1 769 XNOR3X2 $T=2484900 1753360 1 0 $X=2484898 $Y=1747920
X1223 768 6166 776 3 1 7818 XNOR3X2 $T=2523840 1723120 0 0 $X=2523838 $Y=1722718
X1224 7912 7783 7465 3 1 7931 XNOR3X2 $T=2573340 1723120 0 0 $X=2573338 $Y=1722718
X1225 7509 7495 803 3 1 806 XNOR3X2 $T=2594460 1743280 1 0 $X=2594458 $Y=1737840
X1226 796 819 806 3 1 8098 XNOR3X2 $T=2617560 1743280 1 0 $X=2617558 $Y=1737840
X1227 4583 1 401 4586 410 4559 3 AOI22XL $T=1535820 1763440 0 180 $X=1532520 $Y=1758000
X1228 4672 1 430 4633 4640 4641 3 AOI22XL $T=1554300 1642480 0 180 $X=1551000 $Y=1637040
X1229 6767 1 6747 6730 6732 6773 3 AOI22XL $T=2231460 1723120 1 0 $X=2231458 $Y=1717680
X1230 4949 4706 3 1 4572 4931 4947 OAI211X2 $T=1641420 1723120 1 180 $X=1634820 $Y=1722718
X1231 5070 4933 3 1 5050 5007 5072 OAI211X2 $T=1675080 1692880 1 180 $X=1668480 $Y=1692478
X1232 192 89 3 1 BUFX4 $T=1134540 1753360 0 180 $X=1131240 $Y=1747920
X1233 295 95 3 1 BUFX4 $T=1237500 1692880 1 180 $X=1234200 $Y=1692478
X1234 325 200 3 1 BUFX4 $T=1281720 1632400 0 180 $X=1278420 $Y=1626960
X1235 3998 185 3 1 BUFX4 $T=1329240 1763440 1 180 $X=1325940 $Y=1763038
X1236 3928 238 3 1 BUFX4 $T=1336500 1632400 1 180 $X=1333200 $Y=1631998
X1237 401 422 3 1 BUFX4 $T=1535820 1763440 1 0 $X=1535818 $Y=1758000
X1238 5203 483 3 1 BUFX4 $T=1722600 1753360 1 0 $X=1722598 $Y=1747920
X1239 6028 621 3 1 BUFX4 $T=2001120 1753360 1 180 $X=1997820 $Y=1752958
X1240 6015 631 3 1 BUFX4 $T=2018280 1662640 1 0 $X=2018278 $Y=1657200
X1241 4707 4660 3 1 4715 NAND2BX4 $T=1569480 1662640 0 0 $X=1569478 $Y=1662238
X1242 4437 4365 4415 1 3 4419 OR3XL $T=1487640 1723120 0 180 $X=1484340 $Y=1717680
X1243 4432 4365 4415 1 3 4457 OR3XL $T=1486980 1723120 0 0 $X=1486978 $Y=1722718
X1244 4436 4437 3 4438 4432 4403 1 OAI22XL $T=1488300 1733200 0 0 $X=1488298 $Y=1732798
X1245 608 604 3 606 314 611 1 OAI22XL $T=1960860 1763440 1 180 $X=1956900 $Y=1763038
X1246 2538 2536 2510 2515 3 1 AND3X4 $T=903540 1652560 1 180 $X=899580 $Y=1652158
X1247 8054 3 8047 1 8043 7988 NAND3XL $T=2609640 1682800 1 0 $X=2609638 $Y=1677360
X1248 446 444 442 3 4676 1 OAI2BB1XL $T=1584660 1622320 0 180 $X=1581360 $Y=1616880
X1249 7719 7721 7582 3 7730 1 OAI2BB1XL $T=2523180 1763440 0 0 $X=2523178 $Y=1763038
X1250 237 256 3 255 257 1 258 259 250 OAI222X1 $T=1205160 1622320 0 0 $X=1205158 $Y=1621918
X1251 247 256 3 255 203 1 251 259 252 OAI222X1 $T=1207140 1642480 1 0 $X=1207138 $Y=1637040
X1252 243 256 3 255 261 1 240 259 263 OAI222X1 $T=1207800 1652560 1 0 $X=1207798 $Y=1647120
X1253 248 256 3 255 233 1 244 259 264 OAI222X1 $T=1208460 1702960 1 0 $X=1208458 $Y=1697520
X1254 296 256 3 255 282 1 289 259 298 OAI222X1 $T=1249380 1713040 0 0 $X=1249378 $Y=1712638
X1255 293 256 3 255 290 1 323 259 3723 OAI222X1 $T=1294260 1723120 1 0 $X=1294258 $Y=1717680
X1256 332 3 3842 1 CLKINVX8 $T=1315380 1632400 0 0 $X=1315378 $Y=1631998
X1257 433 3 432 1 CLKINVX8 $T=1565520 1713040 1 180 $X=1561560 $Y=1712638
X1258 4765 3 4707 1 CLKINVX8 $T=1587960 1662640 0 0 $X=1587958 $Y=1662238
X1259 4765 3 4685 1 CLKINVX8 $T=1591920 1662640 0 0 $X=1591918 $Y=1662238
X1260 497 3 5303 1 CLKINVX8 $T=1760880 1642480 0 180 $X=1756920 $Y=1637040
X1261 5788 3 598 1 CLKINVX8 $T=1927200 1652560 1 0 $X=1927198 $Y=1647120
X1262 104 193 86 196 194 201 191 3 1 AOI222X4 $T=1146420 1652560 1 180 $X=1138500 $Y=1652158
X1263 3289 3302 1 3 204 NOR2BX4 $T=1141140 1763440 1 0 $X=1141138 $Y=1758000
X1264 4728 4743 4725 1 3 4749 NAND3BX2 $T=1577400 1733200 1 0 $X=1577398 $Y=1727760
X1265 4833 4853 4852 1 3 4400 NAND3BX2 $T=1609740 1672720 1 0 $X=1609738 $Y=1667280
X1266 2478 98 96 3 2478 1 98 96 2477 OAI222XL $T=891000 1743280 0 180 $X=885720 $Y=1737840
X1267 101 83 2509 3 101 1 2509 83 2478 OAI222XL $T=896280 1763440 0 0 $X=896278 $Y=1763038
X1268 2382 2544 104 3 2544 1 2382 104 2575 OAI222XL $T=904200 1713040 0 0 $X=904198 $Y=1712638
X1269 2540 94 2540 3 2542 1 2542 94 2544 OAI222XL $T=904200 1723120 0 0 $X=904198 $Y=1722718
X1270 207 3297 203 3 202 1 200 82 198 OAI222XL $T=1145760 1632400 0 180 $X=1140480 $Y=1626960
X1271 217 216 214 3 212 1 200 92 3134 OAI222XL $T=1176120 1622320 0 180 $X=1170840 $Y=1616880
X1272 217 3448 223 3 202 1 200 2382 3419 OAI222XL $T=1185360 1702960 0 0 $X=1185358 $Y=1702558
X1273 207 2542 233 3 212 1 200 2422 3420 OAI222XL $T=1195260 1733200 0 180 $X=1189980 $Y=1727760
X1274 207 3356 235 3 202 1 200 171 3421 OAI222XL $T=1195920 1753360 0 180 $X=1190640 $Y=1747920
X1275 217 3516 249 3 212 1 200 98 3518 OAI222XL $T=1206480 1753360 0 180 $X=1201200 $Y=1747920
X1276 239 256 255 3 235 1 272 259 3626 OAI222XL $T=1226940 1713040 0 0 $X=1226938 $Y=1712638
X1277 207 2509 282 3 202 1 200 270 3648 OAI222XL $T=1242780 1702960 1 180 $X=1237500 $Y=1702558
X1278 207 2576 261 3 212 1 200 288 280 OAI222XL $T=1238820 1632400 1 0 $X=1238818 $Y=1626960
X1279 207 281 284 3 212 1 200 3651 3612 OAI222XL $T=1240140 1723120 1 0 $X=1240138 $Y=1717680
X1280 217 292 290 3 202 1 200 285 3650 OAI222XL $T=1246080 1753360 0 180 $X=1240800 $Y=1747920
X1281 207 304 305 3 202 1 200 308 3703 OAI222XL $T=1262580 1753360 1 0 $X=1262578 $Y=1747920
X1282 207 139 307 3 212 1 200 3721 3682 OAI222XL $T=1265220 1713040 1 0 $X=1265218 $Y=1707600
X1283 3743 256 255 3 307 1 309 259 3728 OAI222XL $T=1271820 1713040 1 180 $X=1266540 $Y=1712638
X1284 217 318 315 3 212 1 200 313 3775 OAI222XL $T=1287660 1753360 0 180 $X=1282380 $Y=1747920
X1285 302 256 255 3 284 1 333 259 3760 OAI222XL $T=1312740 1723120 1 0 $X=1312738 $Y=1717680
X1286 340 346 255 3 315 1 341 259 3965 OAI222XL $T=1349700 1733200 1 180 $X=1344420 $Y=1732798
X1287 535 514 5463 3 530 1 374 5348 532 OAI222XL $T=1816320 1622320 0 180 $X=1811040 $Y=1616880
X1288 566 550 514 3 557 1 554 538 5555 OAI222XL $T=1846680 1622320 1 180 $X=1841400 $Y=1621918
X1289 5500 550 514 3 561 1 347 538 5559 OAI222XL $T=1847340 1652560 0 180 $X=1842060 $Y=1647120
X1290 548 514 550 3 562 1 214 538 5552 OAI222XL $T=1847340 1692880 1 180 $X=1842060 $Y=1692478
X1291 571 550 514 3 560 1 555 538 5560 OAI222XL $T=1847340 1702960 1 180 $X=1842060 $Y=1702558
X1292 569 5463 514 3 563 1 558 5348 5562 OAI222XL $T=1848000 1672720 1 180 $X=1842720 $Y=1672318
X1293 573 550 514 3 567 1 565 538 570 OAI222XL $T=1849980 1622320 0 180 $X=1844700 $Y=1616880
X1294 3296 3288 3 1 197 AND2X4 $T=1137840 1723120 0 0 $X=1137838 $Y=1722718
X1295 4581 444 3 1 427 AND2X4 $T=1584000 1662640 0 0 $X=1583998 $Y=1662238
X1296 502 503 3 1 5399 AND2X4 $T=1770780 1682800 1 0 $X=1770778 $Y=1677360
X1297 502 455 3 1 5381 AND2X4 $T=1773420 1662640 0 0 $X=1773418 $Y=1662238
X1298 124 120 111 3 1 2728 MX2X1 $T=966900 1773520 0 180 $X=961620 $Y=1768080
X1299 124 122 110 3 1 2731 MX2X1 $T=968220 1662640 1 180 $X=962940 $Y=1662238
X1300 124 123 114 3 1 2732 MX2X1 $T=968220 1692880 1 180 $X=962940 $Y=1692478
X1301 124 130 115 3 1 2756 MX2X1 $T=985380 1723120 0 180 $X=980100 $Y=1717680
X1302 124 157 144 3 1 3000 MX2X1 $T=1050720 1662640 1 180 $X=1045440 $Y=1662238
X1303 3074 1 3 97 BUFX8 $T=1076460 1743280 1 0 $X=1076458 $Y=1737840
X1304 401 1 3 389 BUFX8 $T=1498200 1763440 1 0 $X=1498198 $Y=1758000
X1305 4476 1 3 325 BUFX8 $T=1502820 1622320 1 0 $X=1502818 $Y=1616880
X1306 4769 1 3 4702 BUFX8 $T=1589280 1702960 1 0 $X=1589278 $Y=1697520
X1307 428 1 3 4785 BUFX8 $T=1597860 1713040 0 0 $X=1597858 $Y=1712638
X1308 428 1 3 4798 BUFX8 $T=1599840 1702960 1 0 $X=1599838 $Y=1697520
X1309 410 4529 1 4522 4432 4527 3 AOI22X2 $T=1516680 1753360 1 180 $X=1510740 $Y=1752958
X1310 410 411 1 4522 4457 4510 3 AOI22X2 $T=1518000 1773520 0 180 $X=1512060 $Y=1768080
X1311 4522 4528 1 365 4512 4540 3 AOI22X2 $T=1516020 1733200 0 0 $X=1516018 $Y=1732798
X1312 427 4528 1 4522 425 4616 3 AOI22X2 $T=1554300 1733200 1 180 $X=1548360 $Y=1732798
X1313 4975 4927 1 4949 4917 5006 3 AOI22X2 $T=1655280 1733200 1 180 $X=1649340 $Y=1732798
X1314 506 522 1 5393 518 519 3 AOI22X2 $T=1802460 1682800 1 180 $X=1796520 $Y=1682398
X1315 5381 508 3 1 BUFX16 $T=1787940 1682800 0 0 $X=1787938 $Y=1682398
X1316 5399 509 3 1 BUFX16 $T=1820280 1682800 0 0 $X=1820278 $Y=1682398
X1317 98 97 3 108 1 2591 2604 OAI211XL $T=924660 1773520 0 180 $X=920700 $Y=1768080
X1318 118 117 115 2714 112 1 3 2643 SDFFRHQX1 $T=961620 1763440 0 180 $X=945120 $Y=1758000
X1319 118 117 34 2878 112 1 3 133 SDFFRHQX1 $T=1009140 1763440 0 180 $X=992640 $Y=1758000
X1320 118 117 28 3113 169 1 3 3077 SDFFRHQX1 $T=1086360 1642480 1 180 $X=1069860 $Y=1642078
X1321 118 117 86 3425 169 1 3 3369 SDFFRHQX1 $T=1182060 1702960 0 180 $X=1165560 $Y=1697520
X1322 118 117 185 3895 169 1 3 342 SDFFRHQX1 $T=1319340 1773520 1 0 $X=1319338 $Y=1768080
X1323 364 479 518 5418 483 1 3 5467 SDFFRHQX1 $T=1792560 1672720 1 0 $X=1792558 $Y=1667280
X1324 364 588 5975 5974 491 1 3 5973 SDFFRHQX1 $T=1989900 1713040 1 0 $X=1989898 $Y=1707600
X1325 364 588 633 6056 491 1 3 5975 SDFFRHQX1 $T=2016960 1713040 1 0 $X=2016958 $Y=1707600
X1326 3 1 111 ANTENNA $T=960300 1773520 1 0 $X=960298 $Y=1768080
X1327 3 1 324 ANTENNA $T=1912020 1733200 0 0 $X=1912018 $Y=1732798
X1328 3 1 329 ANTENNA $T=1913340 1723120 0 0 $X=1913338 $Y=1722718
X1329 118 117 30 2780 112 2747 3 1 SDFFRHQX2 $T=988020 1763440 0 180 $X=968220 $Y=1758000
X1330 118 117 139 2867 112 2803 3 1 SDFFRHQX2 $T=1007160 1733200 0 180 $X=987360 $Y=1727760
X1331 118 117 37 3100 169 3074 3 1 SDFFRHQX2 $T=1084380 1733200 0 180 $X=1064580 $Y=1727760
X1332 118 117 97 3109 169 3075 3 1 SDFFRHQX2 $T=1085700 1682800 0 180 $X=1065900 $Y=1677360
X1333 118 117 3651 3650 169 3605 3 1 SDFFRHQX2 $T=1245420 1763440 1 180 $X=1225620 $Y=1763038
X1334 118 117 308 3775 169 327 3 1 SDFFRHQX2 $T=1285020 1773520 1 0 $X=1285018 $Y=1768080
X1335 364 478 501 5334 491 507 3 1 SDFFRHQX2 $T=1762860 1713040 1 0 $X=1762858 $Y=1707600
X1336 364 479 544 532 483 549 3 1 SDFFRHQX2 $T=1828200 1642480 0 0 $X=1828198 $Y=1642078
X1337 364 478 578 5562 491 575 3 1 SDFFRHQX2 $T=1880340 1682800 1 0 $X=1880338 $Y=1677360
X1338 364 588 629 6016 491 620 3 1 SDFFRHQX2 $T=2010360 1773520 0 180 $X=1990560 $Y=1768080
X1339 2747 34 3 1 BUFX12 $T=974820 1763440 0 0 $X=974818 $Y=1763038
X1340 3987 255 3 1 BUFX12 $T=1350360 1713040 1 180 $X=1343760 $Y=1712638
X1341 4015 259 3 1 BUFX12 $T=1365540 1733200 1 180 $X=1358940 $Y=1732798
X1342 5275 487 3 1 BUFX12 $T=1746360 1622320 0 0 $X=1746358 $Y=1621918
X1343 118 88 117 3419 169 1 3 86 SDFFRHQX4 $T=1180740 1692880 0 180 $X=1156320 $Y=1687440
X1344 118 104 117 3420 169 1 3 208 SDFFRHQX4 $T=1180740 1733200 0 180 $X=1156320 $Y=1727760
X1345 118 208 117 3421 169 1 3 192 SDFFRHQX4 $T=1180740 1753360 0 180 $X=1156320 $Y=1747920
X1346 118 210 117 3518 169 1 3 88 SDFFRHQX4 $T=1210440 1763440 0 180 $X=1186020 $Y=1758000
X1347 354 120 117 3965 169 1 3 3998 SDFFRHQX4 $T=1380720 1773520 1 180 $X=1356300 $Y=1773118
X1348 364 489 479 5229 483 1 3 485 SDFFRHQX4 $T=1735140 1642480 0 180 $X=1710720 $Y=1637040
X1349 364 525 478 5478 491 1 3 540 SDFFRHQX4 $T=1806420 1743280 1 0 $X=1806418 $Y=1737840
X1350 364 549 479 5514 483 1 3 518 SDFFRHQX4 $T=1840080 1662640 0 180 $X=1815660 $Y=1657200
X1351 364 577 478 5555 491 1 3 544 SDFFRHQX4 $T=1856580 1632400 1 0 $X=1856578 $Y=1626960
X1352 364 551 478 5559 491 1 3 536 SDFFRHQX4 $T=1859880 1642480 0 0 $X=1859878 $Y=1642078
X1353 364 585 478 5552 491 1 3 578 SDFFRHQX4 $T=1878360 1692880 1 0 $X=1878358 $Y=1687440
X1354 364 520 588 5714 491 1 3 582 SDFFRHQX4 $T=1906080 1773520 1 180 $X=1881660 $Y=1773118
X1355 364 5757 478 5774 491 1 3 585 SDFFRHQX4 $T=1919280 1692880 0 0 $X=1919278 $Y=1692478
X1356 364 543 478 5802 491 1 3 5757 SDFFRHQX4 $T=1950960 1672720 0 180 $X=1926540 $Y=1667280
X1357 3356 219 220 1 215 3450 3 AOI2BB2XL $T=1184040 1713040 0 0 $X=1184038 $Y=1712638
X1358 232 219 221 1 215 3436 3 AOI2BB2XL $T=1189320 1622320 0 180 $X=1184700 $Y=1616880
X1359 3448 219 230 1 215 3461 3 AOI2BB2XL $T=1187340 1682800 0 0 $X=1187338 $Y=1682398
X1360 2542 211 234 1 226 3469 3 AOI2BB2XL $T=1191960 1692880 0 0 $X=1191958 $Y=1692478
X1361 2576 219 236 1 226 3479 3 AOI2BB2XL $T=1193940 1652560 1 0 $X=1193938 $Y=1647120
X1362 2509 3664 287 1 283 3649 3 AOI2BB2XL $T=1244760 1713040 1 180 $X=1240140 $Y=1712638
X1363 139 219 300 1 226 3712 3 AOI2BB2XL $T=1257300 1723120 0 0 $X=1257298 $Y=1722718
X1364 292 219 324 1 283 3819 3 AOI2BB2XL $T=1296240 1733200 0 0 $X=1296238 $Y=1732798
X1365 318 3664 336 1 226 3886 3 AOI2BB2XL $T=1318020 1733200 0 0 $X=1318018 $Y=1732798
X1366 5500 448 503 1 536 5485 3 AOI2BB2XL $T=1821600 1642480 1 180 $X=1816980 $Y=1642078
X1367 227 248 244 238 3469 2714 1 3 OAI221X4 $T=1202520 1702960 0 180 $X=1195260 $Y=1697520
X1368 227 296 289 242 3649 2867 1 3 OAI221X4 $T=1245420 1733200 0 180 $X=1238160 $Y=1727760
X1369 227 3743 309 238 3712 303 1 3 OAI221X4 $T=1273800 1723120 1 180 $X=1266540 $Y=1722718
X1370 227 293 323 242 3819 2878 1 3 OAI221X4 $T=1302840 1733200 0 180 $X=1295580 $Y=1727760
X1371 804 8024 807 801 809 8056 1 3 OAI221X4 $T=2604360 1773520 0 0 $X=2604358 $Y=1773118
X1372 229 256 255 223 260 259 267 1 3 OAI222X4 $T=1206480 1662640 0 0 $X=1206478 $Y=1662238
X1373 265 256 255 249 262 259 254 1 3 OAI222X4 $T=1214400 1713040 1 180 $X=1206480 $Y=1712638
X1374 317 256 255 305 314 259 311 1 3 OAI222X4 $T=1289640 1723120 0 180 $X=1281720 $Y=1717680
X1375 227 265 262 3 238 1 3488 3100 OAI221X1 $T=1213080 1723120 1 180 $X=1207800 $Y=1722718
X1376 8043 7980 7980 3 8047 1 8055 7940 OAI221X1 $T=2606340 1672720 1 0 $X=2606338 $Y=1667280
X1377 118 117 186 3648 169 270 83 3 1 SDFFRX4 $T=1249380 1682800 0 180 $X=1226280 $Y=1677360
X1378 118 117 270 3612 169 3651 295 3 1 SDFFRX4 $T=1226940 1692880 1 0 $X=1226938 $Y=1687440
X1379 118 117 3721 3723 169 293 178 3 1 SDFFRX4 $T=1269180 1652560 0 180 $X=1246080 $Y=1647120
X1380 118 117 278 3682 169 3721 84 3 1 SDFFRX4 $T=1246740 1632400 0 0 $X=1246738 $Y=1631998
X1381 118 117 91 3703 169 308 85 3 1 SDFFRX4 $T=1252020 1773520 1 0 $X=1252018 $Y=1768080
X1382 118 117 184 3760 169 302 186 3 1 SDFFRX4 $T=1283700 1682800 1 180 $X=1260600 $Y=1682398
X1383 3721 3 3651 270 285 3719 1 NAND4X1 $T=1263240 1692880 0 0 $X=1263238 $Y=1692478
X1384 389 1 391 122 3 4327 4351 AOI22X4 $T=1459260 1763440 0 0 $X=1459258 $Y=1763038
X1385 4419 3 4436 4457 1 4438 4275 OAI22X2 $T=1490940 1743280 1 0 $X=1490938 $Y=1737840
X1386 400 3 1 4472 BUFXL $T=1497540 1662640 0 0 $X=1497538 $Y=1662238
X1387 403 3 1 376 BUFXL $T=1506780 1682800 1 0 $X=1506778 $Y=1677360
X1388 4581 3 1 4582 BUFXL $T=1533840 1642480 0 0 $X=1533838 $Y=1642078
X1389 4581 3 1 4590 BUFXL $T=1536480 1652560 1 0 $X=1536478 $Y=1647120
X1390 429 3 1 4672 BUFXL $T=1554960 1632400 1 0 $X=1554958 $Y=1626960
X1391 123 405 4477 1 4400 4325 3 AOI31X2 $T=1500180 1743280 1 0 $X=1500178 $Y=1737840
X1392 5485 527 529 1 526 528 3 AOI31X2 $T=1813020 1652560 0 180 $X=1807080 $Y=1647120
X1393 4513 3 4527 412 1 4327 NAND3X4 $T=1511400 1763440 1 0 $X=1511398 $Y=1758000
X1394 4616 3 4609 4597 1 4397 NAND3X4 $T=1544400 1733200 1 180 $X=1537800 $Y=1732798
X1395 439 3 4716 4742 1 392 NAND3X4 $T=1574100 1713040 0 0 $X=1574098 $Y=1712638
X1396 424 3 4660 426 1 4638 NAND3BX1 $T=1554300 1662640 0 180 $X=1551000 $Y=1657200
X1397 430 3 4837 4831 1 454 NAND3BX1 $T=1605780 1622320 0 180 $X=1602480 $Y=1616880
X1398 4707 3 447 1 4774 4782 410 OAI22X4 $T=1587300 1692880 1 0 $X=1587298 $Y=1687440
X1399 4685 3 447 1 4774 4782 4779 OAI22X4 $T=1589940 1682800 1 0 $X=1589938 $Y=1677360
X1400 428 1 3 4777 BUFX2 $T=1595880 1692880 0 0 $X=1595878 $Y=1692478
X1401 509 1 3 5596 BUFX2 $T=1858560 1682800 0 0 $X=1858558 $Y=1682398
X1402 424 4884 406 4868 3 1 OR3X4 $T=1618320 1652560 1 180 $X=1612380 $Y=1652158
X1403 4885 4849 1 3 4892 4933 NOR3X4 $T=1617660 1702960 1 0 $X=1617658 $Y=1697520
X1404 5005 3 5007 1 CLKINVX2 $T=1650660 1723120 1 0 $X=1650658 $Y=1717680
X1405 5018 3 5014 1 CLKINVX2 $T=1657260 1682800 0 180 $X=1655280 $Y=1677360
X1406 4911 4944 3 5006 457 5036 1 470 OAI221X2 $T=1655280 1753360 0 0 $X=1655278 $Y=1752958
X1407 499 506 3 1 INVX20 $T=1764840 1682800 0 0 $X=1764838 $Y=1682398
X1408 517 494 492 531 1 3 523 NAND4X4 $T=1807080 1702960 0 180 $X=1795860 $Y=1697520
X1409 506 556 1 577 5393 3 5614 581 AOI221X2 $T=1871760 1682800 1 180 $X=1863840 $Y=1682398
X1410 813 8077 1 8080 8020 3 7943 8061 AOI221X2 $T=2620200 1642480 1 180 $X=2612280 $Y=1642078
X1411 5757 5767 5787 1 3 5788 MX2X2 $T=1921260 1652560 1 0 $X=1921258 $Y=1647120
X1412 7864 7777 1 7888 3 7923 7943 AOI211XL $T=2576640 1642480 0 0 $X=2576638 $Y=1642078
X1413 7988 7981 7086 7975 3 1 MXI2X2 $T=2599080 1682800 1 180 $X=2593800 $Y=1682398
.ENDS
***************************************
.SUBCKT CMPR22X1 S A B VDD VSS CO
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB2X2 A0N A1N VSS B1 B0 Y VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDHX1 S A B VDD VSS CO
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX20 A VSS VDD Y
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CMPR42X1 ICO B A C D CO ICI VSS VDD S
** N=12 EP=10 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI31XL A2 A1 VSS A0 B0 Y VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_59 2 3 19 21 22 23 24 27 28 30 31 34 36 37 38 39 40 41 42 43
+ 44 45 46 48 49 50 51 52 53 54 55 57 58 59 61 62 63 64 65 66
+ 67 68 69 70 71 72 73 74 75 77 79 80 81 82 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 125 126 128 129 130 131 133
+ 134 136 137 138 139 140 141 143 144 146 148 149 150 151 152 153 154 155 156 157
+ 158 159 160 161 162 163 164 165 166 167 168 171 172 173 174 176 177 178 179 180
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 223
+ 224 225 226 227 229 230 231 232 233 235 236 238 240 241 242 243 245 246 247 248
+ 249 251 252 253 254 255 257 258 260 262 264 265 266 268 269 270 271 272 273 274
+ 276 277 278 279 281 282 284 286 288 289 291 292 294 296 298 299 300 302 303 304
+ 305 306 307 308 309 310 311 313 314 315 316 317 318 319 320 321 322 323 324 325
+ 326 327 328 329 330 331 333 334 335 337 338 339 340 341 343 345 346 347 348 349
+ 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366 367 368 369
+ 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389
+ 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409
+ 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429
+ 430 431 432 433 435 436 438 439 440 442 443 444 445 446 447 448 449 450 451 452
+ 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472
+ 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492
+ 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512
+ 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530 531 532
+ 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552
+ 553 555 556 557 558 559 561 562 563 564 565 566 567 568 569 571 572 573 574 575
+ 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595
+ 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615
+ 616 618 619 620 621 622 623 624 625 626 627 628 629 631 632 633 634 636 638 639
+ 641 642 644 645 647 648 650 651 652 653 654 656 659 661 662 663 665 666 668 669
+ 670 671 672 673 675 676 677 680 681 683 684 685 686 688 689 690 692 693 694 696
+ 697 699 700 702 705 707 708 709 710 711 713 715 717 718 719 720 721 722 723 724
+ 725 726 727 728 729 730 731 732 736 738 739 741 742 743 744 747 748 749 750 751
+ 752 753 754 755 756 757 758 759 760 761 762 763 764 765 766 767 768 769 770 771
+ 772 773 775 776 777 778 779 780 781 782 783 784 785 786 787 788 789 790 791 792
+ 793 794 795 796 797 798 799 800 801 803 804 806 807 808 809 810 811 812 814 815
+ 817 818 819 820 822 823 824 825 826 827 828 829 830 831 832 833 834 835 836 837
+ 838 839 840 841 842 843 844 845 846 847 848 849 850 851 852 853 858 859 875 1733
+ 1734
** N=31337 EP=741 IP=13307 FDC=0
X0 41 3 42 2 1761 NAND2X1 $T=669240 1914640 0 0 $X=669238 $Y=1914238
X1 1845 3 59 2 1829 NAND2X1 $T=693000 1793680 1 0 $X=692998 $Y=1788240
X2 1963 3 1912 2 66 NAND2X1 $T=716760 1793680 0 0 $X=716758 $Y=1793278
X3 1972 3 1989 2 2050 NAND2X1 $T=727980 1813840 1 180 $X=726000 $Y=1813438
X4 1975 3 1998 2 2049 NAND2X1 $T=735900 1823920 1 0 $X=735898 $Y=1818480
X5 71 3 2052 2 2051 NAND2X1 $T=739860 1965040 1 180 $X=737880 $Y=1964638
X6 77 3 75 2 2136 NAND2X1 $T=750420 1965040 1 180 $X=748440 $Y=1964638
X7 2211 3 2206 2 90 NAND2X1 $T=772860 1783600 0 180 $X=770880 $Y=1778160
X8 2216 3 2275 2 2272 NAND2X1 $T=786720 1975120 1 0 $X=786718 $Y=1969680
X9 2320 3 2363 2 2361 NAND2X1 $T=799920 1803760 1 0 $X=799918 $Y=1798320
X10 2369 3 2367 2 2299 NAND2X1 $T=803880 1844080 1 180 $X=801900 $Y=1843678
X11 2476 3 103 2 2451 NAND2X1 $T=834240 1975120 1 0 $X=834238 $Y=1969680
X12 2469 3 2491 2 2587 NAND2X1 $T=838860 1874320 0 180 $X=836880 $Y=1868880
X13 2587 3 2525 2 2527 NAND2X1 $T=846780 1874320 1 0 $X=846778 $Y=1868880
X14 2586 3 2589 2 2508 NAND2X1 $T=855360 1823920 1 0 $X=855358 $Y=1818480
X15 2613 3 2592 2 2590 NAND2X1 $T=858660 1874320 0 180 $X=856680 $Y=1868880
X16 2591 3 107 2 2517 NAND2X1 $T=857340 1803760 0 0 $X=857338 $Y=1803358
X17 2633 3 2664 2 2638 NAND2X1 $T=873840 1894480 0 0 $X=873838 $Y=1894078
X18 2756 3 2746 2 2820 NAND2X1 $T=894960 1904560 1 180 $X=892980 $Y=1904158
X19 111 3 2753 2 2742 NAND2X1 $T=894300 1834000 1 0 $X=894298 $Y=1828560
X20 2698 3 2700 2 2756 NAND2X1 $T=894300 1914640 0 0 $X=894298 $Y=1914238
X21 109 3 2771 2 2708 NAND2X1 $T=898920 1813840 1 180 $X=896940 $Y=1813438
X22 2773 3 2774 2 2780 NAND2X1 $T=898260 1894480 1 0 $X=898258 $Y=1889040
X23 2772 3 2806 2 2773 NAND2X1 $T=906180 1894480 0 180 $X=904200 $Y=1889040
X24 118 3 2498 2 2878 NAND2X1 $T=922680 1813840 0 180 $X=920700 $Y=1808400
X25 2878 3 2874 2 2895 NAND2X1 $T=925320 1823920 1 0 $X=925318 $Y=1818480
X26 62 3 50 2 2934 NAND2X1 $T=939180 1914640 1 180 $X=937200 $Y=1914238
X27 120 3 2315 2 2939 NAND2X1 $T=942480 1854160 1 0 $X=942478 $Y=1848720
X28 2939 3 2913 2 2948 NAND2X1 $T=942480 1864240 0 0 $X=942478 $Y=1863838
X29 121 3 2317 2 2958 NAND2X1 $T=946440 1793680 1 0 $X=946438 $Y=1788240
X30 2934 3 2935 2 3022 NAND2X1 $T=946440 1924720 1 0 $X=946438 $Y=1919280
X31 2958 3 2917 2 2936 NAND2X1 $T=948420 1803760 0 180 $X=946440 $Y=1798320
X32 68 3 58 2 2947 NAND2X1 $T=947760 1914640 1 0 $X=947758 $Y=1909200
X33 133 3 2840 2 3045 NAND2X1 $T=977460 1854160 1 0 $X=977458 $Y=1848720
X34 2891 3 3114 2 3131 NAND2X1 $T=982740 1884400 0 0 $X=982738 $Y=1883998
X35 3103 3 3106 2 3135 NAND2X1 $T=986700 1904560 0 0 $X=986698 $Y=1904158
X36 3213 3 3142 2 3224 NAND2X1 $T=1004520 1834000 0 180 $X=1002540 $Y=1828560
X37 3212 3 2841 2 3210 NAND2X1 $T=1005180 1864240 1 0 $X=1005178 $Y=1858800
X38 3210 3 3095 2 3258 NAND2X1 $T=1009140 1864240 0 0 $X=1009138 $Y=1863838
X39 150 3 3213 2 3158 NAND2X1 $T=1014420 1834000 0 0 $X=1014418 $Y=1833598
X40 3293 3 3299 2 3311 NAND2X1 $T=1028940 1854160 1 0 $X=1028938 $Y=1848720
X41 3321 3 2842 2 3324 NAND2X1 $T=1035540 1904560 0 0 $X=1035538 $Y=1904158
X42 161 3 163 2 3338 NAND2X1 $T=1043460 1783600 1 0 $X=1043458 $Y=1778160
X43 62 3 111 2 3339 NAND2X1 $T=1044780 1864240 1 0 $X=1044778 $Y=1858800
X44 3457 3 2938 2 3369 NAND2X1 $T=1046100 1894480 1 0 $X=1046098 $Y=1889040
X45 166 3 171 2 3436 NAND2X1 $T=1058640 1894480 1 0 $X=1058638 $Y=1889040
X46 3463 3 3465 2 3435 NAND2X1 $T=1064580 1813840 0 0 $X=1064578 $Y=1813438
X47 3513 3 3514 2 3485 NAND2X1 $T=1075800 1904560 1 0 $X=1075798 $Y=1899120
X48 3485 3 3526 2 3547 NAND2X1 $T=1079760 1914640 1 0 $X=1079758 $Y=1909200
X49 191 3 182 2 3480 NAND2X1 $T=1082400 1783600 1 0 $X=1082398 $Y=1778160
X50 3438 3 3522 2 3574 NAND2X1 $T=1087680 1975120 1 0 $X=1087678 $Y=1969680
X51 190 3 194 2 3582 NAND2X1 $T=1090320 1793680 0 0 $X=1090318 $Y=1793278
X52 3241 3 3592 2 3652 NAND2X1 $T=1094280 1914640 1 0 $X=1094278 $Y=1909200
X53 199 3 198 2 3650 NAND2X1 $T=1103520 1854160 1 0 $X=1103518 $Y=1848720
X54 179 3 187 2 3658 NAND2X1 $T=1103520 1985200 0 0 $X=1103518 $Y=1984798
X55 3659 3 3657 2 3656 NAND2X1 $T=1105500 1894480 0 180 $X=1103520 $Y=1889040
X56 3651 3 3622 2 3659 NAND2X1 $T=1106160 1874320 0 0 $X=1106158 $Y=1873918
X57 205 3 204 2 3674 NAND2X1 $T=1114740 1813840 1 180 $X=1112760 $Y=1813438
X58 55 3 209 2 3813 NAND2X1 $T=1120020 1783600 1 0 $X=1120018 $Y=1778160
X59 53 3 209 2 3760 NAND2X1 $T=1123980 1783600 0 0 $X=1123978 $Y=1783198
X60 3791 3 3152 2 3774 NAND2X1 $T=1136520 1904560 0 180 $X=1134540 $Y=1899120
X61 3878 3 3876 2 3820 NAND2X1 $T=1156980 1884400 1 0 $X=1156978 $Y=1878960
X62 3931 3 3918 2 3913 NAND2X1 $T=1164240 1854160 0 180 $X=1162260 $Y=1848720
X63 3934 3 3058 2 3940 NAND2X1 $T=1166220 1904560 0 0 $X=1166218 $Y=1904158
X64 223 3 3958 2 4118 NAND2X1 $T=1179420 1793680 1 0 $X=1179418 $Y=1788240
X65 4025 3 4033 2 4013 NAND2X1 $T=1189980 1874320 1 0 $X=1189978 $Y=1868880
X66 4079 3 4047 2 3972 NAND2X1 $T=1193940 1864240 1 180 $X=1191960 $Y=1863838
X67 4069 3 220 2 4073 NAND2X1 $T=1197240 1783600 1 0 $X=1197238 $Y=1778160
X68 4145 3 4127 2 4143 NAND2X1 $T=1207140 1904560 0 180 $X=1205160 $Y=1899120
X69 4117 3 3431 2 4145 NAND2X1 $T=1209120 1914640 0 0 $X=1209118 $Y=1914238
X70 4202 3 3460 2 4239 NAND2X1 $T=1226280 1904560 0 0 $X=1226278 $Y=1904158
X71 4235 3 220 2 4255 NAND2X1 $T=1227600 1793680 1 0 $X=1227598 $Y=1788240
X72 112 3 219 2 4283 NAND2X1 $T=1228260 1793680 0 0 $X=1228258 $Y=1793278
X73 4029 3 3789 2 4267 NAND2X1 $T=1230240 1793680 0 0 $X=1230238 $Y=1793278
X74 4277 3 220 2 4281 NAND2X1 $T=1232220 1793680 0 0 $X=1232218 $Y=1793278
X75 115 3 219 2 4238 NAND2X1 $T=1234200 1783600 1 0 $X=1234198 $Y=1778160
X76 4288 3 4312 2 4287 NAND2X1 $T=1242120 1874320 1 0 $X=1242118 $Y=1868880
X77 4358 3 4307 2 4340 NAND2X1 $T=1246740 1965040 0 180 $X=1244760 $Y=1959600
X78 4327 3 3589 2 4304 NAND2X1 $T=1247400 1914640 1 0 $X=1247398 $Y=1909200
X79 4393 3 4395 2 4339 NAND2X1 $T=1252680 1874320 0 0 $X=1252678 $Y=1873918
X80 265 3 264 2 4360 NAND2X1 $T=1259280 1985200 1 180 $X=1257300 $Y=1984798
X81 109 3 219 2 4438 NAND2X1 $T=1257960 1793680 0 0 $X=1257958 $Y=1793278
X82 4410 3 220 2 4430 NAND2X1 $T=1259940 1793680 0 0 $X=1259938 $Y=1793278
X83 4431 3 4396 2 4286 NAND2X1 $T=1261260 1823920 1 0 $X=1261258 $Y=1818480
X84 62 3 3789 2 4437 NAND2X1 $T=1261920 1793680 0 0 $X=1261918 $Y=1793278
X85 4449 3 3932 2 4398 NAND2X1 $T=1264560 1914640 0 180 $X=1262580 $Y=1909200
X86 4407 3 4473 2 4472 NAND2X1 $T=1270500 1944880 1 0 $X=1270498 $Y=1939440
X87 111 3 219 2 4477 NAND2X1 $T=1272480 1793680 1 0 $X=1272478 $Y=1788240
X88 4489 3 4453 2 4417 NAND2X1 $T=1277760 1894480 0 180 $X=1275780 $Y=1889040
X89 4495 3 3010 2 4501 NAND2X1 $T=1278420 1823920 0 0 $X=1278418 $Y=1823518
X90 4503 3 3832 2 4533 NAND2X1 $T=1286340 1904560 0 0 $X=1286338 $Y=1904158
X91 4613 3 4612 2 4632 NAND2X1 $T=1304160 1854160 0 180 $X=1302180 $Y=1848720
X92 286 3 4485 2 4611 NAND2X1 $T=1308780 1874320 1 0 $X=1308778 $Y=1868880
X93 4668 3 3056 2 4693 NAND2X1 $T=1323300 1813840 0 0 $X=1323298 $Y=1813438
X94 4733 3 4694 2 4649 NAND2X1 $T=1327920 1864240 0 180 $X=1325940 $Y=1858800
X95 4766 3 4706 2 4750 NAND2X1 $T=1341780 1844080 1 180 $X=1339800 $Y=1843678
X96 4841 3 4766 2 4779 NAND2X1 $T=1349700 1854160 0 180 $X=1347720 $Y=1848720
X97 321 3 322 2 4880 NAND2X1 $T=1372800 1884400 1 0 $X=1372798 $Y=1878960
X98 326 3 325 2 4930 NAND2X1 $T=1389960 1985200 1 0 $X=1389958 $Y=1979760
X99 334 3 335 2 5081 NAND2X1 $T=1403820 1985200 1 0 $X=1403818 $Y=1979760
X100 5121 3 338 2 5105 NAND2X1 $T=1411080 1793680 1 180 $X=1409100 $Y=1793278
X101 340 3 339 2 5122 NAND2X1 $T=1413720 1985200 1 180 $X=1411740 $Y=1984798
X102 4902 3 5147 2 5161 NAND2X1 $T=1418340 1944880 0 0 $X=1418338 $Y=1944478
X103 5131 3 5161 2 5186 NAND2X1 $T=1422300 1944880 0 180 $X=1420320 $Y=1939440
X104 348 3 5173 2 5213 NAND2X1 $T=1434840 1965040 0 180 $X=1432860 $Y=1959600
X105 5341 3 5252 2 5367 NAND2X1 $T=1463220 1924720 1 0 $X=1463218 $Y=1919280
X106 366 3 5339 2 5321 NAND2X1 $T=1465860 1965040 1 0 $X=1465858 $Y=1959600
X107 374 3 368 2 5385 NAND2X1 $T=1467840 1975120 1 180 $X=1465860 $Y=1974718
X108 379 3 384 2 5442 NAND2X1 $T=1479720 1985200 0 0 $X=1479718 $Y=1984798
X109 5467 3 5523 2 5478 NAND2X1 $T=1495560 1904560 0 0 $X=1495558 $Y=1904158
X110 405 3 401 2 5581 NAND2X1 $T=1513380 1985200 0 180 $X=1511400 $Y=1979760
X111 410 3 407 2 5610 NAND2X1 $T=1519980 1965040 1 180 $X=1518000 $Y=1964638
X112 412 3 5651 2 403 NAND2X1 $T=1524600 1783600 1 0 $X=1524598 $Y=1778160
X113 5651 3 5688 2 5645 NAND2X1 $T=1532520 1793680 1 0 $X=1532518 $Y=1788240
X114 5719 3 402 2 5740 NAND2X1 $T=1539120 1793680 0 180 $X=1537140 $Y=1788240
X115 419 3 409 2 5719 NAND2X1 $T=1540440 1783600 1 0 $X=1540438 $Y=1778160
X116 5746 3 414 2 5695 NAND2X1 $T=1545060 1934800 0 0 $X=1545058 $Y=1934398
X117 421 3 420 2 5724 NAND2X1 $T=1547040 1954960 0 180 $X=1545060 $Y=1949520
X118 5798 3 5799 2 5802 NAND2X1 $T=1552980 1904560 1 0 $X=1552978 $Y=1899120
X119 425 3 409 2 5806 NAND2X1 $T=1555620 1783600 1 0 $X=1555618 $Y=1778160
X120 5804 3 423 2 5836 NAND2X1 $T=1582020 1783600 0 0 $X=1582018 $Y=1783198
X121 5935 3 5912 2 5913 NAND2X1 $T=1584000 1904560 0 180 $X=1582020 $Y=1899120
X122 6014 3 448 2 6061 NAND2X1 $T=1602480 1793680 0 180 $X=1600500 $Y=1788240
X123 6129 3 6080 2 6133 NAND2X1 $T=1638120 1975120 0 180 $X=1636140 $Y=1969680
X124 6239 3 472 2 6222 NAND2X1 $T=1655940 1975120 0 180 $X=1653960 $Y=1969680
X125 6251 3 6256 2 6169 NAND2X1 $T=1663200 1934800 0 0 $X=1663198 $Y=1934398
X126 6299 3 6294 2 6295 NAND2X1 $T=1675740 1924720 0 180 $X=1673760 $Y=1919280
X127 6333 3 479 2 6293 NAND2X1 $T=1675740 1965040 1 180 $X=1673760 $Y=1964638
X128 6377 3 486 2 6299 NAND2X1 $T=1696200 1924720 0 180 $X=1694220 $Y=1919280
X129 6465 3 6449 2 6444 NAND2X1 $T=1708080 1844080 0 180 $X=1706100 $Y=1838640
X130 6451 3 494 2 6501 NAND2X1 $T=1711380 1975120 0 0 $X=1711378 $Y=1974718
X131 6522 3 498 2 6597 NAND2X1 $T=1722600 1894480 1 180 $X=1720620 $Y=1894078
X132 6674 3 507 2 6601 NAND2X1 $T=1742400 1803760 1 180 $X=1740420 $Y=1803358
X133 6699 3 519 2 6673 NAND2X1 $T=1758900 1874320 1 180 $X=1756920 $Y=1873918
X134 6697 3 522 2 6704 NAND2X1 $T=1762860 1793680 0 180 $X=1760880 $Y=1788240
X135 557 3 527 2 6813 NAND2X1 $T=1798500 1844080 1 180 $X=1796520 $Y=1843678
X136 558 3 553 2 6812 NAND2X1 $T=1799820 1975120 1 180 $X=1797840 $Y=1974718
X137 7152 3 7165 2 7167 NAND2X1 $T=1865160 1834000 0 0 $X=1865158 $Y=1833598
X138 520 3 528 2 7152 NAND2X1 $T=1867800 1834000 1 0 $X=1867798 $Y=1828560
X139 7189 3 601 2 7187 NAND2X1 $T=1869780 1934800 0 180 $X=1867800 $Y=1929360
X140 603 3 527 2 7165 NAND2X1 $T=1871760 1834000 0 0 $X=1871758 $Y=1833598
X141 7367 3 7372 2 7384 NAND2X1 $T=1937760 1944880 1 0 $X=1937758 $Y=1939440
X142 611 3 7407 2 7472 NAND2X1 $T=1937760 1944880 0 0 $X=1937758 $Y=1944478
X143 625 3 7543 2 7525 NAND2X1 $T=1963500 1934800 0 180 $X=1961520 $Y=1929360
X144 473 3 7609 2 7615 NAND2X1 $T=1978020 1834000 1 0 $X=1978018 $Y=1828560
X145 629 3 7657 2 7646 NAND2X1 $T=1987260 1904560 0 0 $X=1987258 $Y=1904158
X146 633 3 632 2 631 NAND2X1 $T=1989240 1985200 1 180 $X=1987260 $Y=1984798
X147 7616 3 7643 2 7698 NAND2X1 $T=1997820 1965040 1 0 $X=1997818 $Y=1959600
X148 7679 3 7699 2 7660 NAND2X1 $T=1998480 1944880 0 0 $X=1998478 $Y=1944478
X149 636 3 7683 2 7570 NAND2X1 $T=2001780 1884400 1 0 $X=2001778 $Y=1878960
X150 7782 3 7762 2 7745 NAND2X1 $T=2014980 1844080 0 0 $X=2014978 $Y=1843678
X151 7779 3 7822 2 7866 NAND2X1 $T=2024220 1975120 0 0 $X=2024218 $Y=1974718
X152 644 3 648 2 7799 NAND2X1 $T=2034120 1864240 0 0 $X=2034118 $Y=1863838
X153 7879 3 7840 2 651 NAND2X1 $T=2036100 1965040 1 180 $X=2034120 $Y=1964638
X154 651 3 7866 2 7883 NAND2X1 $T=2038080 1975120 1 180 $X=2036100 $Y=1974718
X155 7878 3 650 2 7818 NAND2X1 $T=2036760 1803760 1 0 $X=2036758 $Y=1798320
X156 653 3 654 2 7856 NAND2X1 $T=2042040 1884400 1 0 $X=2042038 $Y=1878960
X157 7547 3 663 2 7974 NAND2X1 $T=2068440 1783600 1 0 $X=2068438 $Y=1778160
X158 7881 3 8039 2 673 NAND2X1 $T=2077680 1975120 1 0 $X=2077678 $Y=1969680
X159 672 3 669 2 8056 NAND2X1 $T=2086260 1884400 0 0 $X=2086258 $Y=1883998
X160 676 3 625 2 8089 NAND2X1 $T=2094840 1783600 0 0 $X=2094838 $Y=1783198
X161 680 3 681 2 8169 NAND2X1 $T=2103420 1874320 0 180 $X=2101440 $Y=1868880
X162 8052 3 8091 2 8110 NAND2X1 $T=2102100 1965040 1 0 $X=2102098 $Y=1959600
X163 8117 3 8189 2 8184 NAND2X1 $T=2104740 1985200 1 0 $X=2104738 $Y=1979760
X164 684 3 685 2 8170 NAND2X1 $T=2109360 1834000 1 0 $X=2109358 $Y=1828560
X165 8096 3 8212 2 8233 NAND2X1 $T=2116620 1944880 0 0 $X=2116618 $Y=1944478
X166 7098 3 607 2 8257 NAND2X1 $T=2123220 1884400 1 0 $X=2123218 $Y=1878960
X167 8211 3 8273 2 696 NAND2X1 $T=2136420 1944880 1 0 $X=2136418 $Y=1939440
X168 8310 3 8288 2 8316 NAND2X1 $T=2140380 1954960 1 0 $X=2140378 $Y=1949520
X169 8315 3 8365 2 710 NAND2X1 $T=2162820 1975120 0 0 $X=2162818 $Y=1974718
X170 7234 3 541 2 8492 NAND2X1 $T=2183280 1884400 1 0 $X=2183278 $Y=1878960
X171 8496 3 708 2 8527 NAND2X1 $T=2186580 1823920 0 180 $X=2184600 $Y=1818480
X172 8397 3 8495 2 8505 NAND2X1 $T=2189880 1944880 1 0 $X=2189878 $Y=1939440
X173 8512 3 8541 2 8595 NAND2X1 $T=2195160 1965040 1 0 $X=2195158 $Y=1959600
X174 8619 3 8624 2 8660 NAND2X1 $T=2212320 1975120 0 0 $X=2212318 $Y=1974718
X175 8582 3 8584 2 8639 NAND2X1 $T=2216280 1944880 0 0 $X=2216278 $Y=1944478
X176 8599 3 8798 2 8887 NAND2X1 $T=2281620 1944880 1 0 $X=2281618 $Y=1939440
X177 8889 3 8783 2 8978 NAND2X1 $T=2284260 1894480 1 0 $X=2284258 $Y=1889040
X178 8920 3 8921 2 742 NAND2X1 $T=2292840 1975120 0 180 $X=2290860 $Y=1969680
X179 8800 3 8776 2 8993 NAND2X1 $T=2296140 1854160 0 0 $X=2296138 $Y=1853758
X180 8939 3 8780 2 8977 NAND2X1 $T=2297460 1834000 0 0 $X=2297458 $Y=1833598
X181 8831 3 8779 2 9028 NAND2X1 $T=2301420 1834000 1 0 $X=2301418 $Y=1828560
X182 8777 3 8814 2 9041 NAND2X1 $T=2306700 1954960 1 0 $X=2306698 $Y=1949520
X183 9031 3 9023 2 8995 NAND2X1 $T=2313300 1844080 1 180 $X=2311320 $Y=1843678
X184 8797 3 8833 2 9069 NAND2X1 $T=2311980 1914640 1 0 $X=2311978 $Y=1909200
X185 9028 3 9031 2 9033 NAND2X1 $T=2313300 1834000 1 0 $X=2313298 $Y=1828560
X186 9045 3 748 2 751 NAND2X1 $T=2315940 1985200 1 180 $X=2313960 $Y=1984798
X187 8795 3 8832 2 9072 NAND2X1 $T=2316600 1924720 0 0 $X=2316598 $Y=1924318
X188 8812 3 9042 2 9045 NAND2X1 $T=2319240 1975120 1 0 $X=2319238 $Y=1969680
X189 8977 3 9023 2 9111 NAND2X1 $T=2325840 1844080 1 0 $X=2325838 $Y=1838640
X190 9137 3 9120 2 8904 NAND2X1 $T=2334420 1823920 0 180 $X=2332440 $Y=1818480
X191 9121 3 9113 2 9130 NAND2X1 $T=2335080 1924720 0 0 $X=2335078 $Y=1924318
X192 9142 3 9156 2 9094 NAND2X1 $T=2340360 1965040 1 0 $X=2340358 $Y=1959600
X193 9167 3 758 2 9052 NAND2X1 $T=2348280 1803760 1 0 $X=2348278 $Y=1798320
X194 8978 3 9109 2 9227 NAND2X1 $T=2350920 1894480 0 0 $X=2350918 $Y=1894078
X195 9023 3 9240 2 9163 NAND2X1 $T=2358840 1854160 1 0 $X=2358838 $Y=1848720
X196 9241 3 9269 2 9245 NAND2X1 $T=2360160 1965040 0 0 $X=2360158 $Y=1964638
X197 9109 3 9026 2 9298 NAND2X1 $T=2361480 1894480 0 0 $X=2361478 $Y=1894078
X198 9270 3 9317 2 9307 NAND2X1 $T=2377320 1924720 1 0 $X=2377318 $Y=1919280
X199 9316 3 9318 2 9320 NAND2X1 $T=2377320 1965040 1 0 $X=2377318 $Y=1959600
X200 9346 3 9242 2 9321 NAND2X1 $T=2379300 1975120 1 180 $X=2377320 $Y=1974718
X201 9457 3 9456 2 9454 NAND2X1 $T=2402400 1924720 1 180 $X=2400420 $Y=1924318
X202 9458 3 9472 2 9473 NAND2X1 $T=2404380 1884400 0 0 $X=2404378 $Y=1883998
X203 9477 3 9492 2 9455 NAND2X1 $T=2406360 1904560 1 0 $X=2406358 $Y=1899120
X204 9497 3 9500 2 9504 NAND2X1 $T=2412300 1844080 1 0 $X=2412298 $Y=1838640
X205 9274 3 9576 2 9550 NAND2X1 $T=2428140 1904560 1 0 $X=2428138 $Y=1899120
X206 9599 3 9627 2 9518 NAND2X1 $T=2440020 1975120 0 0 $X=2440018 $Y=1974718
X207 790 3 9741 2 9726 NAND2X1 $T=2459820 1985200 1 0 $X=2459818 $Y=1979760
X208 9741 3 791 2 9795 NAND2X1 $T=2475660 1985200 0 0 $X=2475658 $Y=1984798
X209 9759 3 9811 2 9814 NAND2X1 $T=2480280 1844080 1 0 $X=2480278 $Y=1838640
X210 9922 3 791 2 9920 NAND2X1 $T=2500080 1965040 0 180 $X=2498100 $Y=1959600
X211 808 3 9944 2 9924 NAND2X1 $T=2511300 1944880 1 180 $X=2509320 $Y=1944478
X212 10088 3 819 2 10053 NAND2X1 $T=2533080 1934800 0 180 $X=2531100 $Y=1929360
X213 827 3 826 2 10227 NAND2X1 $T=2549580 1793680 1 0 $X=2549578 $Y=1788240
X214 10248 3 830 2 10253 NAND2X1 $T=2562780 1954960 1 0 $X=2562778 $Y=1949520
X215 10216 3 828 2 10269 NAND2X1 $T=2564760 1813840 0 0 $X=2564758 $Y=1813438
X216 10253 3 10268 2 10228 NAND2X1 $T=2568060 1914640 1 0 $X=2568058 $Y=1909200
X217 10303 3 836 2 10233 NAND2X1 $T=2580600 1944880 0 180 $X=2578620 $Y=1939440
X218 850 3 849 2 10360 NAND2X1 $T=2609640 1985200 0 0 $X=2609638 $Y=1984798
X219 390 2 3 126 5527 NOR2X4 $T=1495560 1844080 0 0 $X=1495558 $Y=1843678
X220 5527 2 3 5586 5557 NOR2X4 $T=1508100 1844080 0 0 $X=1508098 $Y=1843678
X221 6660 2 3 6659 515 NOR2X4 $T=1754940 1965040 1 0 $X=1754938 $Y=1959600
X222 6678 2 3 6695 488 NOR2X4 $T=1762860 1965040 1 0 $X=1762858 $Y=1959600
X223 1814 3 1829 61 2 NAND2BX1 $T=689700 1783600 0 0 $X=689698 $Y=1783198
X224 2063 3 2051 2090 2 NAND2BX1 $T=743160 1934800 0 0 $X=743158 $Y=1934398
X225 2086 3 2136 2194 2 NAND2BX1 $T=759000 1934800 1 0 $X=758998 $Y=1929360
X226 2294 3 2299 2282 2 NAND2BX1 $T=794640 1844080 1 180 $X=792000 $Y=1843678
X227 2297 3 2361 2381 2 NAND2BX1 $T=799260 1813840 0 0 $X=799258 $Y=1813438
X228 2492 3 2508 2511 2 NAND2BX1 $T=841500 1834000 1 0 $X=841498 $Y=1828560
X229 2490 3 2517 2479 2 NAND2BX1 $T=846780 1823920 1 180 $X=844140 $Y=1823518
X230 2617 3 2590 2709 2 NAND2BX1 $T=877800 1874320 1 0 $X=877798 $Y=1868880
X231 2729 3 2708 2703 2 NAND2BX1 $T=885720 1834000 1 180 $X=883080 $Y=1833598
X232 2754 3 2742 2805 2 NAND2BX1 $T=904200 1844080 0 0 $X=904198 $Y=1843678
X233 3115 3 3131 3138 2 NAND2BX1 $T=985380 1894480 1 0 $X=985378 $Y=1889040
X234 3096 3 3135 3211 2 NAND2BX1 $T=995940 1904560 0 0 $X=995938 $Y=1904158
X235 109 3 152 3163 2 NAND2BX1 $T=1016400 1813840 1 180 $X=1013760 $Y=1813438
X236 3294 3 3311 3417 2 NAND2BX1 $T=1040160 1864240 0 0 $X=1040158 $Y=1863838
X237 3359 3 3369 3437 2 NAND2BX1 $T=1046760 1904560 1 0 $X=1046758 $Y=1899120
X238 3620 3 3582 3566 2 NAND2BX1 $T=1092300 1803760 1 180 $X=1089660 $Y=1803358
X239 3655 3 3652 3711 2 NAND2BX1 $T=1109460 1914640 1 0 $X=1109458 $Y=1909200
X240 3879 3 3774 3893 2 NAND2BX1 $T=1152360 1904560 1 0 $X=1152358 $Y=1899120
X241 3944 3 3940 3917 2 NAND2BX1 $T=1170840 1904560 0 0 $X=1170838 $Y=1904158
X242 4008 3 4003 4034 2 NAND2BX1 $T=1189320 1914640 1 0 $X=1189318 $Y=1909200
X243 4226 3 4239 4264 2 NAND2BX1 $T=1233540 1904560 0 0 $X=1233538 $Y=1904158
X244 249 3 4231 4347 2 NAND2BX1 $T=1238160 1944880 1 0 $X=1238158 $Y=1939440
X245 4411 3 4398 4436 2 NAND2BX1 $T=1259940 1904560 0 0 $X=1259938 $Y=1904158
X246 296 3 294 4562 2 NAND2BX1 $T=1316040 1985200 1 180 $X=1313400 $Y=1984798
X247 4653 3 4673 4672 2 NAND2BX1 $T=1322640 1884400 0 180 $X=1320000 $Y=1878960
X248 4929 3 4789 4923 2 NAND2BX1 $T=1374780 1844080 0 180 $X=1372140 $Y=1838640
X249 4985 3 4967 4914 2 NAND2BX1 $T=1385340 1944880 0 180 $X=1382700 $Y=1939440
X250 5079 3 5081 5010 2 NAND2BX1 $T=1403820 1924720 0 180 $X=1401180 $Y=1919280
X251 5084 3 5104 5168 2 NAND2BX1 $T=1420980 1854160 1 0 $X=1420978 $Y=1848720
X252 5217 3 5202 5188 2 NAND2BX1 $T=1432860 1924720 0 180 $X=1430220 $Y=1919280
X253 5368 3 5385 5359 2 NAND2BX1 $T=1467840 1934800 1 180 $X=1465200 $Y=1934398
X254 5474 3 5438 5477 2 NAND2BX1 $T=1487640 1944880 1 0 $X=1487638 $Y=1939440
X255 5692 3 5695 5700 2 NAND2BX1 $T=1534500 1924720 0 0 $X=1534498 $Y=1924318
X256 5715 3 5724 5713 2 NAND2BX1 $T=1545060 1894480 1 180 $X=1542420 $Y=1894078
X257 5806 3 5651 5804 2 NAND2BX1 $T=1563540 1783600 1 0 $X=1563538 $Y=1778160
X258 433 3 5651 5883 2 NAND2BX1 $T=1566180 1793680 1 0 $X=1566178 $Y=1788240
X259 5838 3 5862 5877 2 NAND2BX1 $T=1571460 1884400 0 0 $X=1571458 $Y=1883998
X260 6291 3 6276 6221 2 NAND2BX1 $T=1670460 1914640 0 180 $X=1667820 $Y=1909200
X261 6447 3 6450 6401 2 NAND2BX1 $T=1704780 1944880 1 180 $X=1702140 $Y=1944478
X262 6446 3 6448 6400 2 NAND2BX1 $T=1714680 1934800 0 180 $X=1712040 $Y=1929360
X263 517 3 516 6660 2 NAND2BX1 $T=1772760 1944880 0 0 $X=1772758 $Y=1944478
X264 603 3 7173 615 2 NAND2BX1 $T=1895520 1975120 0 0 $X=1895518 $Y=1974718
X265 603 3 7173 7235 2 NAND2BX1 $T=1896840 1965040 1 0 $X=1896838 $Y=1959600
X266 7620 3 7570 7571 2 NAND2BX1 $T=1971420 1884400 0 180 $X=1968780 $Y=1878960
X267 7613 3 7615 7589 2 NAND2BX1 $T=1980660 1834000 1 180 $X=1978020 $Y=1833598
X268 7744 3 7745 7676 2 NAND2BX1 $T=2005080 1854160 1 180 $X=2002440 $Y=1853758
X269 7862 3 7856 7816 2 NAND2BX1 $T=2034120 1884400 0 180 $X=2031480 $Y=1878960
X270 625 3 626 7837 2 NAND2BX1 $T=2032800 1823920 0 0 $X=2032798 $Y=1823518
X271 7926 3 7929 7924 2 NAND2BX1 $T=2051280 1783600 1 180 $X=2048640 $Y=1783198
X272 7978 3 7974 7975 2 NAND2BX1 $T=2057880 1803760 0 180 $X=2055240 $Y=1798320
X273 8054 3 8056 8002 2 NAND2BX1 $T=2080980 1894480 0 180 $X=2078340 $Y=1889040
X274 8107 3 8110 677 2 NAND2BX1 $T=2094180 1975120 1 0 $X=2094178 $Y=1969680
X275 8182 3 8170 8111 2 NAND2BX1 $T=2106060 1834000 0 180 $X=2103420 $Y=1828560
X276 9068 3 9069 9304 2 NAND2BX1 $T=2321880 1914640 1 0 $X=2321878 $Y=1909200
X277 754 3 9094 753 2 NAND2BX1 $T=2331120 1985200 0 180 $X=2328480 $Y=1979760
X278 9527 3 9456 9520 2 NAND2BX1 $T=2418900 1965040 0 180 $X=2416260 $Y=1959600
X279 10231 3 10253 10263 2 NAND2BX1 $T=2564760 1904560 0 0 $X=2564758 $Y=1904158
X280 834 3 838 10327 2 NAND2BX1 $T=2579280 1985200 0 0 $X=2579278 $Y=1984798
X281 832 3 841 10429 2 NAND2BX1 $T=2604360 1944880 1 0 $X=2604358 $Y=1939440
X282 66 1814 3 1829 2 1932 OAI21X1 $T=712140 1783600 0 180 $X=708840 $Y=1778160
X283 205 3712 3 3716 2 3564 OAI21X1 $T=1116720 1954960 0 0 $X=1116718 $Y=1954558
X284 4008 4045 3 4003 2 3993 OAI21X1 $T=1182720 1904560 1 180 $X=1179420 $Y=1904158
X285 7744 7677 3 7745 2 7761 OAI21X1 $T=1998480 1844080 0 0 $X=1998478 $Y=1843678
X286 7819 7862 3 7856 2 7853 OAI21X1 $T=2034780 1874320 1 180 $X=2031480 $Y=1873918
X287 7998 639 3 7547 2 8038 OAI21X1 $T=2079000 1793680 1 180 $X=2075700 $Y=1793278
X288 7902 8184 3 8218 2 8254 OAI21X1 $T=2112000 1985200 1 0 $X=2111998 $Y=1979760
X289 8308 705 3 8395 2 8396 OAI21X1 $T=2157540 1783600 1 180 $X=2154240 $Y=1783198
X290 9480 9454 3 9483 2 9378 OAI21X1 $T=2405700 1934800 0 0 $X=2405698 $Y=1934398
X291 9527 9505 3 9480 2 785 OAI21X1 $T=2428140 1965040 1 180 $X=2424840 $Y=1964638
X292 2492 3 2477 2508 2 2478 OAI21XL $T=838860 1834000 0 180 $X=836220 $Y=1828560
X293 2508 3 2490 2517 2 2446 OAI21XL $T=844140 1813840 1 180 $X=841500 $Y=1813438
X294 2590 3 2488 2587 2 2588 OAI21XL $T=857340 1874320 1 180 $X=854700 $Y=1873918
X295 2617 3 2656 2590 2 2653 OAI21XL $T=872520 1874320 0 180 $X=869880 $Y=1868880
X296 2742 3 2729 2708 2 2727 OAI21XL $T=891000 1834000 0 180 $X=888360 $Y=1828560
X297 2773 3 2702 2756 2 2693 OAI21XL $T=897600 1894480 1 180 $X=894960 $Y=1894078
X298 2754 3 2781 2742 2 2724 OAI21XL $T=901560 1844080 1 180 $X=898920 $Y=1843678
X299 3135 3 3115 3131 2 3064 OAI21XL $T=988020 1904560 0 180 $X=985380 $Y=1899120
X300 3096 3 3174 3135 2 3225 OAI21XL $T=997260 1904560 1 0 $X=997258 $Y=1899120
X301 3339 3 3294 3311 2 3121 OAI21XL $T=1029600 1864240 1 180 $X=1026960 $Y=1863838
X302 3359 3 3366 3369 2 3322 OAI21XL $T=1046100 1904560 0 0 $X=1046098 $Y=1904158
X303 3515 3 3465 3463 2 3429 OAI21XL $T=1067220 1803760 0 180 $X=1064580 $Y=1798320
X304 3477 3 3438 3522 2 3543 OAI21XL $T=1077120 1965040 0 0 $X=1077118 $Y=1964638
X305 3620 3 3567 3582 2 3479 OAI21XL $T=1100220 1793680 1 180 $X=1097580 $Y=1793278
X306 3673 3 3655 3652 2 3495 OAI21XL $T=1104180 1914640 0 180 $X=1101540 $Y=1909200
X307 50 3 150 3790 2 3794 OAI21XL $T=1140480 1793680 1 0 $X=1140478 $Y=1788240
X308 3879 3 3892 3774 2 3914 OAI21XL $T=1157640 1904560 1 0 $X=1157638 $Y=1899120
X309 3774 3 3944 3940 2 3963 OAI21XL $T=1168200 1904560 1 0 $X=1168198 $Y=1899120
X310 4226 3 4224 4239 2 4125 OAI21XL $T=1223640 1904560 0 180 $X=1221000 $Y=1899120
X311 4366 3 4364 4339 2 4261 OAI21XL $T=1252020 1864240 0 180 $X=1249380 $Y=1858800
X312 4408 3 4411 4398 2 4313 OAI21XL $T=1257300 1904560 1 180 $X=1254660 $Y=1904158
X313 4520 3 4527 4516 2 4440 OAI21XL $T=1285020 1864240 1 180 $X=1282380 $Y=1863838
X314 4632 3 4650 4649 2 4636 OAI21XL $T=1312080 1854160 0 0 $X=1312078 $Y=1853758
X315 4611 3 4653 4673 2 4486 OAI21XL $T=1316040 1884400 1 180 $X=1313400 $Y=1883998
X316 4930 3 4985 4967 2 4999 OAI21XL $T=1389300 1944880 1 0 $X=1389298 $Y=1939440
X317 5079 3 5078 5081 2 5030 OAI21XL $T=1401840 1934800 0 180 $X=1399200 $Y=1929360
X318 5081 3 5089 5122 2 5108 OAI21XL $T=1409100 1965040 1 0 $X=1409098 $Y=1959600
X319 5212 3 5210 5213 2 5204 OAI21XL $T=1434840 1904560 1 180 $X=1432200 $Y=1904158
X320 5213 3 5217 5202 2 5228 OAI21XL $T=1434840 1934800 1 0 $X=1434838 $Y=1929360
X321 5367 3 5210 5426 2 5424 OAI21XL $T=1477080 1914640 1 0 $X=1477078 $Y=1909200
X322 5442 3 5474 5438 2 5428 OAI21XL $T=1482360 1944880 0 180 $X=1479720 $Y=1939440
X323 5582 3 5426 5569 2 5565 OAI21XL $T=1506780 1924720 1 180 $X=1504140 $Y=1924318
X324 5581 3 5609 5610 2 5566 OAI21XL $T=1513380 1954960 1 0 $X=1513378 $Y=1949520
X325 5612 3 5559 5581 2 5606 OAI21XL $T=1516020 1914640 1 180 $X=1513380 $Y=1914238
X326 5210 3 5633 5629 2 5632 OAI21XL $T=1518660 1904560 1 0 $X=1518658 $Y=1899120
X327 5715 3 5568 5724 2 5696 OAI21XL $T=1538460 1894480 1 180 $X=1535820 $Y=1894078
X328 5724 3 5692 5695 2 5743 OAI21XL $T=1543740 1924720 0 0 $X=1543738 $Y=1924318
X329 5802 3 5568 5800 2 5771 OAI21XL $T=1559580 1874320 1 180 $X=1556940 $Y=1873918
X330 5837 3 5800 5841 2 5844 OAI21XL $T=1563540 1884400 1 0 $X=1563538 $Y=1878960
X331 5913 3 5568 5902 2 5901 OAI21XL $T=1584000 1914640 0 180 $X=1581360 $Y=1909200
X332 6215 3 6291 6276 2 6292 OAI21XL $T=1681020 1914640 1 0 $X=1681018 $Y=1909200
X333 6399 3 6446 6448 2 493 OAI21XL $T=1701480 1934800 1 0 $X=1701478 $Y=1929360
X334 6349 3 6447 6450 2 6482 OAI21XL $T=1710060 1954960 1 0 $X=1710058 $Y=1949520
X335 6815 3 6862 6861 2 6877 OAI21XL $T=1802460 1803760 1 0 $X=1802458 $Y=1798320
X336 6798 3 6753 6800 2 6920 OAI21XL $T=1803780 1813840 0 0 $X=1803778 $Y=1813438
X337 6806 3 550 6810 2 6862 OAI21XL $T=1807080 1793680 1 0 $X=1807078 $Y=1788240
X338 6892 3 557 6893 2 6960 OAI21XL $T=1819620 1844080 0 0 $X=1819618 $Y=1843678
X339 6961 3 6960 6922 2 6982 OAI21XL $T=1828200 1844080 0 0 $X=1828198 $Y=1843678
X340 7566 3 7613 7615 2 7618 OAI21XL $T=1978020 1844080 0 0 $X=1978018 $Y=1843678
X341 7586 3 7620 7570 2 7636 OAI21XL $T=1980000 1884400 1 0 $X=1979998 $Y=1878960
X342 7851 3 647 7854 2 645 OAI21XL $T=2031480 1985200 1 180 $X=2028840 $Y=1984798
X343 7974 3 7926 7929 2 7977 OAI21XL $T=2060520 1783600 0 180 $X=2057880 $Y=1778160
X344 673 3 8107 8110 2 8130 OAI21XL $T=2102100 1975120 1 0 $X=2102098 $Y=1969680
X345 8213 3 689 8232 2 8090 OAI21XL $T=2115960 1783600 1 0 $X=2115958 $Y=1778160
X346 696 3 8314 8316 2 8312 OAI21XL $T=2138400 1965040 0 0 $X=2138398 $Y=1964638
X347 8308 3 8272 689 2 8232 OAI21XL $T=2141040 1783600 0 180 $X=2138400 $Y=1778160
X348 8445 3 7547 8473 2 8496 OAI21XL $T=2180640 1803760 1 0 $X=2180638 $Y=1798320
X349 710 3 8504 8505 2 8602 OAI21XL $T=2187240 1975120 0 0 $X=2187238 $Y=1974718
X350 8532 3 8511 8527 2 8526 OAI21XL $T=2195160 1823920 1 180 $X=2192520 $Y=1823518
X351 8595 3 8600 8639 2 8623 OAI21XL $T=2218260 1965040 0 180 $X=2215620 $Y=1959600
X352 8978 3 8905 8919 2 9021 OAI21XL $T=2299440 1884400 0 0 $X=2299438 $Y=1883998
X353 8887 3 9032 9041 2 9040 OAI21XL $T=2317260 1944880 0 180 $X=2314620 $Y=1939440
X354 9072 3 9068 9069 2 9112 OAI21XL $T=2324520 1924720 1 0 $X=2324518 $Y=1919280
X355 8983 3 9090 8993 2 9075 OAI21XL $T=2329800 1854160 1 180 $X=2327160 $Y=1853758
X356 8992 3 9114 8887 2 9108 OAI21XL $T=2333100 1944880 1 180 $X=2330460 $Y=1944478
X357 761 3 9239 760 2 9162 OAI21XL $T=2358840 1783600 1 0 $X=2358838 $Y=1778160
X358 765 3 9239 9279 2 9280 OAI21XL $T=2368740 1803760 0 0 $X=2368738 $Y=1803358
X359 9114 3 9298 9164 2 9286 OAI21XL $T=2374020 1894480 0 180 $X=2371380 $Y=1889040
X360 768 3 9325 764 2 9356 OAI21XL $T=2383260 1793680 1 0 $X=2383258 $Y=1788240
X361 9520 3 9505 9517 2 9460 OAI21XL $T=2417580 1965040 1 180 $X=2414940 $Y=1964638
X362 9484 3 781 780 2 9525 OAI21XL $T=2420220 1793680 1 180 $X=2417580 $Y=1793278
X363 9538 3 9568 9486 2 9571 OAI21XL $T=2430120 1864240 0 180 $X=2427480 $Y=1858800
X364 786 3 9722 9543 2 9723 OAI21XL $T=2460480 1844080 0 180 $X=2457840 $Y=1838640
X365 787 3 788 9724 2 9744 OAI21XL $T=2464440 1783600 0 0 $X=2464438 $Y=1783198
X366 793 3 789 9744 2 9745 OAI21XL $T=2464440 1813840 1 0 $X=2464438 $Y=1808400
X367 800 3 797 798 2 9837 OAI21XL $T=2492820 1783600 0 180 $X=2490180 $Y=1778160
X368 806 3 9872 808 2 10003 OAI21XL $T=2508660 1965040 0 0 $X=2508658 $Y=1964638
X369 812 3 9964 810 2 9963 OAI21XL $T=2512620 1813840 1 180 $X=2509980 $Y=1813438
X370 804 3 9971 9963 2 9976 OAI21XL $T=2512620 1834000 1 0 $X=2512618 $Y=1828560
X371 823 3 817 820 2 10152 OAI21XL $T=2546940 1803760 0 180 $X=2544300 $Y=1798320
X372 2278 94 2317 3 2 XOR2X4 $T=787380 1783600 0 0 $X=787378 $Y=1783198
X373 2936 2964 3056 3 2 XOR2X4 $T=941820 1813840 1 0 $X=941818 $Y=1808400
X374 8982 8937 744 3 2 XOR2X4 $T=2305380 1813840 0 180 $X=2294160 $Y=1808400
X375 796 9778 795 3 2 XOR2X4 $T=2480280 1975120 0 180 $X=2469060 $Y=1969680
X376 9924 9868 801 3 2 XOR2X4 $T=2505360 1934800 0 180 $X=2494140 $Y=1929360
X377 10054 10032 814 3 2 XOR2X4 $T=2532420 1904560 1 180 $X=2521200 $Y=1904158
X378 10327 10318 835 3 2 XOR2X4 $T=2589180 1894480 0 180 $X=2577960 $Y=1889040
X379 10429 10406 844 3 2 XOR2X4 $T=2607000 1934800 1 180 $X=2595780 $Y=1934398
X380 851 10410 846 3 2 XOR2X4 $T=2608320 1965040 1 180 $X=2597100 $Y=1964638
X381 2086 3 2 2067 INVX1 $T=746460 1934800 0 180 $X=745140 $Y=1929360
X382 2050 3 2 2138 INVX1 $T=758340 1813840 1 0 $X=758338 $Y=1808400
X383 82 3 2 2250 INVX1 $T=764280 1813840 0 180 $X=762960 $Y=1808400
X384 2272 3 2 2274 INVX1 $T=791340 1944880 0 180 $X=790020 $Y=1939440
X385 2364 3 2 2279 INVX1 $T=802560 1944880 1 0 $X=802558 $Y=1939440
X386 2294 3 2 2401 INVX1 $T=821040 1834000 1 0 $X=821038 $Y=1828560
X387 2477 3 2 2447 INVX1 $T=832920 1834000 0 180 $X=831600 $Y=1828560
X388 106 3 2 2500 INVX1 $T=842160 1783600 0 0 $X=842158 $Y=1783198
X389 2488 3 2 2525 INVX1 $T=844800 1884400 1 0 $X=844798 $Y=1878960
X390 2526 3 2 2477 INVX1 $T=848100 1834000 1 180 $X=846780 $Y=1833598
X391 2702 3 2 2746 INVX1 $T=877140 1904560 1 180 $X=875820 $Y=1904158
X392 2731 3 2 2774 INVX1 $T=887700 1884400 1 180 $X=886380 $Y=1883998
X393 114 3 2 2753 INVX1 $T=894300 1793680 0 0 $X=894298 $Y=1793278
X394 115 3 2 2771 INVX1 $T=896940 1783600 1 0 $X=896938 $Y=1778160
X395 2773 3 2 2807 INVX1 $T=907500 1894480 0 0 $X=907498 $Y=1894078
X396 2660 3 2 2697 INVX1 $T=913440 1894480 0 0 $X=913438 $Y=1894078
X397 2749 3 2 2781 INVX1 $T=919380 1844080 0 180 $X=918060 $Y=1838640
X398 2899 3 2 2900 INVX1 $T=926640 1823920 1 180 $X=925320 $Y=1823518
X399 2934 3 2 2930 INVX1 $T=940500 1924720 0 180 $X=939180 $Y=1919280
X400 2939 3 2 2902 INVX1 $T=942480 1854160 1 180 $X=941160 $Y=1853758
X401 2947 3 2 2933 INVX1 $T=943140 1924720 1 180 $X=941820 $Y=1924318
X402 2958 3 2 2932 INVX1 $T=947760 1793680 1 180 $X=946440 $Y=1793278
X403 3045 3 2 3062 INVX1 $T=962280 1854160 0 0 $X=962278 $Y=1853758
X404 3163 3 2 3142 INVX1 $T=996600 1823920 0 0 $X=996598 $Y=1823518
X405 3121 3 2 3174 INVX1 $T=999240 1894480 1 0 $X=999238 $Y=1889040
X406 3210 3 2 3067 INVX1 $T=1000560 1864240 0 180 $X=999240 $Y=1858800
X407 112 3 2 3213 INVX1 $T=1015740 1834000 0 180 $X=1014420 $Y=1828560
X408 3324 3 2 3295 INVX1 $T=1031580 1914640 1 180 $X=1030260 $Y=1914238
X409 156 3 2 158 INVX1 $T=1032900 1783600 1 0 $X=1032898 $Y=1778160
X410 168 3 2 166 INVX1 $T=1047420 1934800 0 180 $X=1046100 $Y=1929360
X411 3357 3 2 3458 INVX1 $T=1061940 1934800 0 0 $X=1061938 $Y=1934398
X412 3485 3 2 3484 INVX1 $T=1069860 1914640 0 0 $X=1069858 $Y=1914238
X413 174 3 2 160 INVX1 $T=1080420 1944880 1 0 $X=1080418 $Y=1939440
X414 3564 3 2 3521 INVX1 $T=1083720 1884400 0 180 $X=1082400 $Y=1878960
X415 3650 3 2 3610 INVX1 $T=1102200 1844080 0 180 $X=1100880 $Y=1838640
X416 3659 3 2 3698 INVX1 $T=1108800 1884400 1 0 $X=1108798 $Y=1878960
X417 3674 3 2 3609 INVX1 $T=1110120 1823920 1 180 $X=1108800 $Y=1823518
X418 3715 3 2 3689 INVX1 $T=1118040 1904560 0 180 $X=1116720 $Y=1899120
X419 176 3 2 192 INVX1 $T=1129260 1803760 1 0 $X=1129258 $Y=1798320
X420 3897 3 2 3749 INVX1 $T=1149720 1854160 1 180 $X=1148400 $Y=1853758
X421 3993 3 2 3892 INVX1 $T=1157640 1894480 1 180 $X=1156320 $Y=1894078
X422 3913 3 2 3939 INVX1 $T=1160940 1834000 0 0 $X=1160938 $Y=1833598
X423 50 3 2 215 INVX1 $T=1176780 1783600 0 0 $X=1176778 $Y=1783198
X424 4013 3 2 3985 INVX1 $T=1183380 1874320 0 180 $X=1182060 $Y=1868880
X425 4145 3 2 4122 INVX1 $T=1207800 1914640 0 180 $X=1206480 $Y=1909200
X426 58 3 2 251 INVX1 $T=1231560 1823920 0 0 $X=1231558 $Y=1823518
X427 246 3 2 4231 INVX1 $T=1232880 1944880 1 0 $X=1232878 $Y=1939440
X428 4340 3 2 4199 INVX1 $T=1234200 1944880 1 180 $X=1232880 $Y=1944478
X429 4287 3 2 4251 INVX1 $T=1235520 1864240 0 180 $X=1234200 $Y=1858800
X430 4304 3 2 4310 INVX1 $T=1238820 1914640 1 0 $X=1238818 $Y=1909200
X431 257 3 2 4358 INVX1 $T=1249380 1965040 1 180 $X=1248060 $Y=1964638
X432 4417 3 2 4432 INVX1 $T=1260600 1874320 0 0 $X=1260598 $Y=1873918
X433 4407 3 2 4456 INVX1 $T=1263240 1934800 0 0 $X=1263238 $Y=1934398
X434 3991 3 2 4470 INVX1 $T=1273800 1813840 0 0 $X=1273798 $Y=1813438
X435 4533 3 2 4480 INVX1 $T=1283040 1904560 0 180 $X=1281720 $Y=1899120
X436 4501 3 2 4555 INVX1 $T=1289640 1823920 1 0 $X=1289638 $Y=1818480
X437 4636 3 2 4520 INVX1 $T=1298220 1854160 1 180 $X=1296900 $Y=1853758
X438 4693 3 2 4629 INVX1 $T=1316700 1803760 1 180 $X=1315380 $Y=1803358
X439 4472 3 2 4706 INVX1 $T=1320660 1844080 0 0 $X=1320658 $Y=1843678
X440 68 3 2 281 INVX1 $T=1321980 1783600 1 180 $X=1320660 $Y=1783198
X441 4842 3 2 4841 INVX1 $T=1356300 1854160 0 180 $X=1354980 $Y=1848720
X442 318 3 2 4902 INVX1 $T=1362900 1954960 1 0 $X=1362898 $Y=1949520
X443 4789 3 2 4917 INVX1 $T=1370160 1834000 0 0 $X=1370158 $Y=1833598
X444 4971 3 2 4915 INVX1 $T=1371480 1954960 1 180 $X=1370160 $Y=1954558
X445 4921 3 2 4928 INVX1 $T=1381380 1834000 1 0 $X=1381378 $Y=1828560
X446 4863 3 2 5025 INVX1 $T=1397880 1793680 1 180 $X=1396560 $Y=1793278
X447 4923 3 2 5027 INVX1 $T=1403160 1844080 1 180 $X=1401840 $Y=1843678
X448 5079 3 2 5102 INVX1 $T=1405140 1924720 0 0 $X=1405138 $Y=1924318
X449 4999 3 2 5078 INVX1 $T=1409760 1924720 0 0 $X=1409758 $Y=1924318
X450 5165 3 2 5167 INVX1 $T=1422960 1803760 1 0 $X=1422958 $Y=1798320
X451 5228 3 2 5258 INVX1 $T=1436160 1924720 0 0 $X=1436158 $Y=1924318
X452 5235 3 2 352 INVX1 $T=1439460 1854160 1 180 $X=1438140 $Y=1853758
X453 333 3 2 360 INVX1 $T=1461900 1783600 0 0 $X=1461898 $Y=1783198
X454 5387 3 2 5396 INVX1 $T=1467180 1854160 1 0 $X=1467178 $Y=1848720
X455 5385 3 2 5399 INVX1 $T=1467180 1944880 0 0 $X=1467178 $Y=1944478
X456 5403 3 2 5368 INVX1 $T=1475100 1965040 0 180 $X=1473780 $Y=1959600
X457 367 3 2 5383 INVX1 $T=1485000 1823920 1 0 $X=1484998 $Y=1818480
X458 5473 3 2 5445 INVX1 $T=1488300 1934800 1 0 $X=1488298 $Y=1929360
X459 5447 3 2 5499 INVX1 $T=1488960 1783600 1 0 $X=1488958 $Y=1778160
X460 5367 3 2 5523 INVX1 $T=1490940 1914640 0 0 $X=1490938 $Y=1914238
X461 5428 3 2 5559 INVX1 $T=1501500 1934800 0 0 $X=1501498 $Y=1934398
X462 5564 3 2 5582 INVX1 $T=1507440 1934800 1 180 $X=1506120 $Y=1934398
X463 5426 3 2 5605 INVX1 $T=1511400 1904560 1 0 $X=1511398 $Y=1899120
X464 403 3 2 5603 INVX1 $T=1512720 1783600 0 180 $X=1511400 $Y=1778160
X465 5645 3 2 5611 INVX1 $T=1518660 1793680 0 180 $X=1517340 $Y=1788240
X466 5612 3 2 5589 INVX1 $T=1527240 1924720 1 0 $X=1527238 $Y=1919280
X467 5719 3 2 5688 INVX1 $T=1539120 1783600 1 180 $X=1537800 $Y=1783198
X468 433 3 2 5796 INVX1 $T=1564860 1793680 0 180 $X=1563540 $Y=1788240
X469 5863 3 2 5835 INVX1 $T=1570800 1793680 0 0 $X=1570798 $Y=1793278
X470 5844 3 2 5861 INVX1 $T=1572120 1884400 1 0 $X=1572118 $Y=1878960
X471 5883 3 2 5860 INVX1 $T=1576080 1793680 1 180 $X=1574760 $Y=1793278
X472 442 3 2 5967 INVX1 $T=1589940 1834000 0 0 $X=1589938 $Y=1833598
X473 148 3 2 454 INVX1 $T=1613700 1803760 0 0 $X=1613698 $Y=1803358
X474 123 3 2 6143 INVX1 $T=1637460 1854160 0 0 $X=1637458 $Y=1853758
X475 6152 3 2 6215 INVX1 $T=1646040 1914640 0 0 $X=1646038 $Y=1914238
X476 6169 3 2 6218 INVX1 $T=1647360 1944880 1 0 $X=1647358 $Y=1939440
X477 6222 3 2 6135 INVX1 $T=1656600 1965040 0 180 $X=1655280 $Y=1959600
X478 6293 3 2 6321 INVX1 $T=1686960 1965040 1 0 $X=1686958 $Y=1959600
X479 6299 3 2 6361 INVX1 $T=1693560 1914640 1 180 $X=1692240 $Y=1914238
X480 238 3 2 354 INVX1 $T=1723260 1985200 1 0 $X=1723258 $Y=1979760
X481 6501 3 2 6540 INVX1 $T=1729860 1975120 0 0 $X=1729858 $Y=1974718
X482 6660 3 2 6599 INVX1 $T=1749660 1954960 1 180 $X=1748340 $Y=1954558
X483 531 3 2 6723 INVX1 $T=1774740 1834000 0 180 $X=1773420 $Y=1828560
X484 500 3 2 6789 INVX1 $T=1781340 1813840 0 0 $X=1781338 $Y=1813438
X485 512 3 2 6787 INVX1 $T=1783980 1793680 1 0 $X=1783978 $Y=1788240
X486 503 3 2 6798 INVX1 $T=1783980 1803760 0 0 $X=1783978 $Y=1803358
X487 523 3 2 6806 INVX1 $T=1791240 1783600 0 0 $X=1791238 $Y=1783198
X488 6812 3 2 6821 INVX1 $T=1804440 1985200 0 0 $X=1804438 $Y=1984798
X489 501 3 2 6863 INVX1 $T=1807080 1834000 0 0 $X=1807078 $Y=1833598
X490 509 3 2 6892 INVX1 $T=1807080 1854160 1 0 $X=1807078 $Y=1848720
X491 579 3 2 580 INVX1 $T=1825560 1813840 0 180 $X=1824240 $Y=1808400
X492 496 3 2 7014 INVX1 $T=1828200 1834000 0 0 $X=1828198 $Y=1833598
X493 6926 3 2 6936 INVX1 $T=1838760 1975120 0 0 $X=1838758 $Y=1974718
X494 574 3 2 6999 INVX1 $T=1842720 1834000 0 180 $X=1841400 $Y=1828560
X495 7097 3 2 7123 INVX1 $T=1854600 1854160 1 0 $X=1854598 $Y=1848720
X496 7173 3 2 6239 INVX1 $T=1865820 1975120 0 180 $X=1864500 $Y=1969680
X497 520 3 2 7172 INVX1 $T=1867140 1823920 1 0 $X=1867138 $Y=1818480
X498 610 3 2 7147 INVX1 $T=1881660 1823920 1 180 $X=1880340 $Y=1823518
X499 7245 3 2 473 INVX1 $T=1892880 1823920 0 180 $X=1891560 $Y=1818480
X500 559 3 2 7173 INVX1 $T=1895520 1975120 0 180 $X=1894200 $Y=1969680
X501 7384 3 2 7421 INVX1 $T=1929840 1975120 1 0 $X=1929838 $Y=1969680
X502 616 3 2 7245 INVX1 $T=1933800 1823920 1 0 $X=1933798 $Y=1818480
X503 7350 3 2 7425 INVX1 $T=1937760 1844080 0 0 $X=1937758 $Y=1843678
X504 626 3 2 7367 INVX1 $T=1960200 1844080 0 180 $X=1958880 $Y=1838640
X505 7525 3 2 7542 INVX1 $T=1961520 1965040 0 0 $X=1961518 $Y=1964638
X506 559 3 2 7407 INVX1 $T=1970100 1944880 0 0 $X=1970098 $Y=1944478
X507 7610 3 2 7639 INVX1 $T=1977360 1975120 1 0 $X=1977358 $Y=1969680
X508 7618 3 2 7677 INVX1 $T=1987920 1844080 0 0 $X=1987918 $Y=1843678
X509 7646 3 2 7587 INVX1 $T=1989240 1894480 1 180 $X=1987920 $Y=1894078
X510 7660 3 2 7662 INVX1 $T=1989240 1965040 1 0 $X=1989238 $Y=1959600
X511 7781 3 2 7609 INVX1 $T=2014980 1823920 1 180 $X=2013660 $Y=1823518
X512 7799 3 2 7813 INVX1 $T=2016300 1874320 1 0 $X=2016298 $Y=1868880
X513 603 3 2 7305 INVX1 $T=2019600 1924720 0 180 $X=2018280 $Y=1919280
X514 7818 3 2 7820 INVX1 $T=2024220 1803760 0 0 $X=2024218 $Y=1803358
X515 7779 3 2 7854 INVX1 $T=2029500 1975120 1 0 $X=2029498 $Y=1969680
X516 7861 3 2 7862 INVX1 $T=2033460 1894480 0 180 $X=2032140 $Y=1889040
X517 7852 3 2 7926 INVX1 $T=2034780 1783600 1 0 $X=2034778 $Y=1778160
X518 7864 3 2 7878 INVX1 $T=2034780 1793680 0 0 $X=2034778 $Y=1793278
X519 656 3 2 7822 INVX1 $T=2047980 1975120 0 0 $X=2047978 $Y=1974718
X520 7961 3 2 7782 INVX1 $T=2054580 1844080 0 180 $X=2053260 $Y=1838640
X521 7978 3 2 7995 INVX1 $T=2062500 1803760 0 180 $X=2061180 $Y=1798320
X522 8006 3 2 7982 INVX1 $T=2067780 1874320 0 180 $X=2066460 $Y=1868880
X523 7960 3 2 7981 INVX1 $T=2068440 1823920 1 0 $X=2068438 $Y=1818480
X524 7902 3 2 665 INVX1 $T=2071740 1985200 1 180 $X=2070420 $Y=1984798
X525 8075 3 2 671 INVX1 $T=2085600 1985200 1 180 $X=2084280 $Y=1984798
X526 8233 3 2 8217 INVX1 $T=2114640 1965040 1 180 $X=2113320 $Y=1964638
X527 8169 3 2 8187 INVX1 $T=2123880 1854160 0 0 $X=2123878 $Y=1853758
X528 550 3 2 7129 INVX1 $T=2126520 1844080 0 0 $X=2126518 $Y=1843678
X529 8254 3 2 694 INVX1 $T=2129160 1985200 0 0 $X=2129158 $Y=1984798
X530 8257 3 2 8412 INVX1 $T=2141700 1884400 1 0 $X=2141698 $Y=1878960
X531 8272 3 2 8395 INVX1 $T=2152260 1783600 1 0 $X=2152258 $Y=1778160
X532 8492 3 2 8539 INVX1 $T=2189220 1884400 1 0 $X=2189218 $Y=1878960
X533 8625 3 2 8530 INVX1 $T=2220240 1813840 1 0 $X=2220238 $Y=1808400
X534 8602 3 2 8782 INVX1 $T=2246640 1975120 0 0 $X=2246638 $Y=1974718
X535 8596 3 2 8679 INVX1 $T=2250600 1975120 0 180 $X=2249280 $Y=1969680
X536 8796 3 2 8835 INVX1 $T=2267760 1985200 1 0 $X=2267758 $Y=1979760
X537 748 3 2 8981 INVX1 $T=2308020 1985200 0 180 $X=2306700 $Y=1979760
X538 9031 3 2 9029 INVX1 $T=2315280 1844080 0 0 $X=2315278 $Y=1843678
X539 9052 3 2 9018 INVX1 $T=2317920 1793680 0 0 $X=2317918 $Y=1793278
X540 9021 3 2 9090 INVX1 $T=2325180 1864240 1 0 $X=2325178 $Y=1858800
X541 8996 3 2 9109 INVX1 $T=2330460 1894480 0 0 $X=2330458 $Y=1894078
X542 9130 3 2 9026 INVX1 $T=2337720 1904560 0 0 $X=2337718 $Y=1904158
X543 9000 3 2 9138 INVX1 $T=2338380 1884400 1 0 $X=2338378 $Y=1878960
X544 8983 3 2 9240 INVX1 $T=2348280 1854160 0 0 $X=2348278 $Y=1853758
X545 9026 3 2 9221 INVX1 $T=2348940 1874320 0 0 $X=2348938 $Y=1873918
X546 9191 3 2 9223 INVX1 $T=2358180 1874320 0 180 $X=2356860 $Y=1868880
X547 9237 3 2 9235 INVX1 $T=2357520 1944880 0 0 $X=2357518 $Y=1944478
X548 8622 3 2 9239 INVX1 $T=2358840 1813840 1 0 $X=2358838 $Y=1808400
X549 9245 3 2 9287 INVX1 $T=2369400 1975120 0 0 $X=2369398 $Y=1974718
X550 768 3 2 9279 INVX1 $T=2377320 1793680 0 0 $X=2377318 $Y=1793278
X551 771 3 2 9325 INVX1 $T=2381280 1783600 1 180 $X=2379960 $Y=1783198
X552 764 3 2 9363 INVX1 $T=2393160 1813840 1 0 $X=2393158 $Y=1808400
X553 9320 3 2 9371 INVX1 $T=2395800 1975120 1 0 $X=2395798 $Y=1969680
X554 9455 3 2 9475 INVX1 $T=2400420 1954960 1 0 $X=2400418 $Y=1949520
X555 9473 3 2 9479 INVX1 $T=2406360 1914640 0 0 $X=2406358 $Y=1914238
X556 778 3 2 9500 INVX1 $T=2409000 1823920 1 0 $X=2408998 $Y=1818480
X557 9550 3 2 9551 INVX1 $T=2421540 1934800 1 0 $X=2421538 $Y=1929360
X558 9480 3 2 9540 INVX1 $T=2424180 1954960 0 180 $X=2422860 $Y=1949520
X559 9568 3 2 9494 INVX1 $T=2426820 1854160 0 0 $X=2426818 $Y=1853758
X560 9538 3 2 9629 INVX1 $T=2442660 1854160 1 0 $X=2442658 $Y=1848720
X561 9599 3 2 9589 INVX1 $T=2442660 1934800 0 0 $X=2442658 $Y=1934398
X562 9593 3 2 9634 INVX1 $T=2442660 1944880 0 0 $X=2442658 $Y=1944478
X563 9627 3 2 9594 INVX1 $T=2443320 1975120 0 0 $X=2443318 $Y=1974718
X564 9706 3 2 9722 INVX1 $T=2458500 1834000 0 0 $X=2458498 $Y=1833598
X565 792 3 2 9741 INVX1 $T=2463120 1985200 0 0 $X=2463118 $Y=1984798
X566 9761 3 2 9762 INVX1 $T=2469060 1864240 0 0 $X=2469058 $Y=1863838
X567 9814 3 2 9835 INVX1 $T=2497440 1864240 1 0 $X=2497438 $Y=1858800
X568 803 3 2 9872 INVX1 $T=2502720 1975120 0 0 $X=2502718 $Y=1974718
X569 804 3 2 9964 INVX1 $T=2510640 1803760 0 0 $X=2510638 $Y=1803358
X570 9836 3 2 9999 INVX1 $T=2510640 1864240 0 0 $X=2510638 $Y=1863838
X571 806 3 2 9944 INVX1 $T=2511960 1954960 0 180 $X=2510640 $Y=1949520
X572 9831 3 2 9972 INVX1 $T=2513280 1874320 0 0 $X=2513278 $Y=1873918
X573 812 3 2 9971 INVX1 $T=2518560 1834000 1 0 $X=2518558 $Y=1828560
X574 10064 3 2 9977 INVX1 $T=2534400 1864240 1 0 $X=2534398 $Y=1858800
X575 10127 3 2 10088 INVX1 $T=2541000 1944880 0 180 $X=2539680 $Y=1939440
X576 10083 3 2 10090 INVX1 $T=2544960 1844080 0 0 $X=2544958 $Y=1843678
X577 10227 3 2 10266 INVX1 $T=2558160 1793680 0 0 $X=2558158 $Y=1793278
X578 10148 3 2 10248 INVX1 $T=2560800 1965040 1 0 $X=2560798 $Y=1959600
X579 832 3 2 10321 INVX1 $T=2573340 1944880 0 0 $X=2573338 $Y=1944478
X580 10233 3 2 10286 INVX1 $T=2577300 1914640 1 180 $X=2575980 $Y=1914238
X581 10254 3 2 10290 INVX1 $T=2589180 1914640 0 0 $X=2589178 $Y=1914238
X582 847 3 2 10412 INVX1 $T=2599740 1783600 0 0 $X=2599738 $Y=1783198
X583 850 3 2 10413 INVX1 $T=2603700 1985200 1 180 $X=2602380 $Y=1984798
X584 845 3 2 10431 INVX1 $T=2608980 1783600 1 180 $X=2607660 $Y=1783198
X585 875 3 2 853 INVX1 $T=2629440 1793680 1 0 $X=2629438 $Y=1788240
X586 1974 69 2 1932 1993 3 AOI21X2 $T=723360 1783600 1 180 $X=718740 $Y=1783198
X587 2900 2874 2 2911 2964 3 AOI21X2 $T=930600 1823920 1 0 $X=930598 $Y=1818480
X588 2911 2917 2 2932 2910 3 AOI21X2 $T=936540 1803760 1 0 $X=936538 $Y=1798320
X589 3810 3880 2 3939 3962 3 AOI21X2 $T=1164900 1823920 0 0 $X=1164898 $Y=1823518
X590 3986 3993 2 3963 3991 3 AOI21X2 $T=1181400 1904560 0 180 $X=1176780 $Y=1899120
X591 7853 7976 2 7982 8004 3 AOI21X2 $T=2056560 1874320 0 0 $X=2056558 $Y=1873918
X592 8051 8119 2 8187 8115 3 AOI21X2 $T=2104740 1854160 0 0 $X=2104738 $Y=1853758
X593 8254 8307 2 8312 8317 3 AOI21X2 $T=2135760 1975120 0 0 $X=2135758 $Y=1974718
X594 9593 9589 2 9551 9480 3 AOI21X2 $T=2432100 1934800 1 180 $X=2427480 $Y=1934398
X595 9966 791 2 10003 10009 3 AOI21X2 $T=2515920 1965040 1 0 $X=2515918 $Y=1959600
X596 10219 10056 2 10228 10032 3 AOI21X2 $T=2556180 1914640 1 0 $X=2556178 $Y=1909200
X597 10303 837 2 833 10254 3 AOI21X2 $T=2580600 1954960 1 180 $X=2575980 $Y=1954558
X598 10056 10325 2 10320 10318 3 AOI21X2 $T=2585880 1934800 1 180 $X=2581260 $Y=1934398
X599 10056 836 2 837 10406 3 AOI21X2 $T=2601060 1954960 0 180 $X=2596440 $Y=1949520
X600 2 1972 1989 1997 3 NOR2X1 $T=727980 1823920 1 180 $X=726000 $Y=1823518
X601 2 2211 2206 89 3 NOR2X1 $T=774180 1783600 1 0 $X=774178 $Y=1778160
X602 2 2369 2367 2294 3 NOR2X1 $T=803220 1834000 0 0 $X=803218 $Y=1833598
X603 2 101 2383 2455 3 NOR2X1 $T=826980 1975120 1 0 $X=826978 $Y=1969680
X604 2 2480 2455 2471 3 NOR2X1 $T=835560 1965040 0 180 $X=833580 $Y=1959600
X605 2 2476 103 2480 3 NOR2X1 $T=836220 1975120 1 180 $X=834240 $Y=1974718
X606 2 2492 2490 2450 3 NOR2X1 $T=838200 1823920 1 180 $X=836220 $Y=1823518
X607 2 2591 107 2490 3 NOR2X1 $T=850740 1803760 1 180 $X=848760 $Y=1803358
X608 2 2586 2589 2492 3 NOR2X1 $T=857340 1834000 0 180 $X=855360 $Y=1828560
X609 2 2488 2617 2633 3 NOR2X1 $T=864600 1884400 0 180 $X=862620 $Y=1878960
X610 2 2613 2592 2617 3 NOR2X1 $T=864600 1874320 1 0 $X=864598 $Y=1868880
X611 2 2614 2499 2639 3 NOR2X1 $T=868560 1965040 0 180 $X=866580 $Y=1959600
X612 2 113 2636 2666 3 NOR2X1 $T=877800 1823920 1 180 $X=875820 $Y=1823518
X613 2 2698 2700 2702 3 NOR2X1 $T=882420 1914640 1 0 $X=882418 $Y=1909200
X614 2 2702 2731 2664 3 NOR2X1 $T=891000 1894480 1 180 $X=889020 $Y=1894078
X615 2 2729 2754 2730 3 NOR2X1 $T=896280 1844080 0 180 $X=894300 $Y=1838640
X616 2 109 2771 2729 3 NOR2X1 $T=898920 1823920 1 180 $X=896940 $Y=1823518
X617 2 111 2753 2754 3 NOR2X1 $T=906180 1834000 1 180 $X=904200 $Y=1833598
X618 2 2772 2806 2731 3 NOR2X1 $T=909480 1884400 0 180 $X=907500 $Y=1878960
X619 2 68 2818 2858 3 NOR2X1 $T=918720 1934800 0 0 $X=918718 $Y=1934398
X620 2 3115 3096 3069 3 NOR2X1 $T=976800 1904560 0 180 $X=974820 $Y=1899120
X621 2 3103 3106 3096 3 NOR2X1 $T=979440 1904560 0 0 $X=979438 $Y=1904158
X622 2 2891 3114 3115 3 NOR2X1 $T=980100 1894480 0 0 $X=980098 $Y=1894078
X623 2 3163 3158 2749 3 NOR2X1 $T=994620 1844080 0 180 $X=992640 $Y=1838640
X624 2 3293 3299 3294 3 NOR2X1 $T=1028940 1854160 0 0 $X=1028938 $Y=1853758
X625 2 3457 2938 3359 3 NOR2X1 $T=1040820 1894480 1 0 $X=1040818 $Y=1889040
X626 2 3241 3592 3655 3 NOR2X1 $T=1096920 1904560 1 0 $X=1096918 $Y=1899120
X627 2 190 194 3620 3 NOR2X1 $T=1108140 1793680 1 180 $X=1106160 $Y=1793278
X628 2 3791 3152 3879 3 NOR2X1 $T=1139820 1904560 1 0 $X=1139818 $Y=1899120
X629 2 3878 3876 3873 3 NOR2X1 $T=1151040 1884400 0 180 $X=1149060 $Y=1878960
X630 2 3934 3058 3944 3 NOR2X1 $T=1162260 1904560 1 180 $X=1160280 $Y=1904158
X631 2 3879 3944 3986 3 NOR2X1 $T=1172160 1904560 1 0 $X=1172158 $Y=1899120
X632 2 4030 3475 4008 3 NOR2X1 $T=1184040 1914640 1 180 $X=1182060 $Y=1914238
X633 2 4178 4126 4128 3 NOR2X1 $T=1213740 1874320 1 180 $X=1211760 $Y=1873918
X634 2 4202 3460 4226 3 NOR2X1 $T=1218360 1914640 1 0 $X=1218358 $Y=1909200
X635 2 4340 4347 4407 3 NOR2X1 $T=1246080 1944880 1 0 $X=1246078 $Y=1939440
X636 2 260 4360 4307 3 NOR2X1 $T=1254660 1985200 0 180 $X=1252680 $Y=1979760
X637 2 4431 4396 4311 3 NOR2X1 $T=1255980 1823920 0 180 $X=1254000 $Y=1818480
X638 2 4393 4395 4364 3 NOR2X1 $T=1255320 1884400 0 0 $X=1255318 $Y=1883998
X639 2 4449 3932 4411 3 NOR2X1 $T=1267200 1904560 1 180 $X=1265220 $Y=1904158
X640 2 276 279 4473 3 NOR2X1 $T=1281720 1944880 0 180 $X=1279740 $Y=1939440
X641 2 4550 4532 4527 3 NOR2X1 $T=1288980 1884400 0 180 $X=1287000 $Y=1878960
X642 2 4562 282 265 3 NOR2X1 $T=1294920 1985200 1 180 $X=1292940 $Y=1984798
X643 2 4684 3933 4653 3 NOR2X1 $T=1325940 1884400 0 0 $X=1325938 $Y=1883998
X644 2 4733 4694 4650 3 NOR2X1 $T=1335180 1864240 0 180 $X=1333200 $Y=1858800
X645 2 304 299 4766 3 NOR2X1 $T=1342440 1864240 1 0 $X=1342438 $Y=1858800
X646 2 4472 4779 4789 3 NOR2X1 $T=1346400 1844080 0 0 $X=1346398 $Y=1843678
X647 2 4921 4917 4920 3 NOR2X1 $T=1372140 1834000 0 180 $X=1370160 $Y=1828560
X648 2 326 325 4971 3 NOR2X1 $T=1384020 1985200 0 180 $X=1382040 $Y=1979760
X649 2 4985 4971 4998 3 NOR2X1 $T=1386000 1954960 1 0 $X=1385998 $Y=1949520
X650 2 328 327 4985 3 NOR2X1 $T=1391940 1954960 1 180 $X=1389960 $Y=1954558
X651 2 334 335 5079 3 NOR2X1 $T=1402500 1975120 1 0 $X=1402498 $Y=1969680
X652 2 5079 5089 5106 3 NOR2X1 $T=1403820 1954960 0 0 $X=1403818 $Y=1954558
X653 2 5028 5088 5104 3 NOR2X1 $T=1409100 1854160 1 0 $X=1409098 $Y=1848720
X654 2 340 339 5089 3 NOR2X1 $T=1419000 1985200 0 0 $X=1418998 $Y=1984798
X655 2 348 5173 5212 3 NOR2X1 $T=1435500 1965040 1 0 $X=1435498 $Y=1959600
X656 2 5199 5236 5217 3 NOR2X1 $T=1441440 1944880 0 180 $X=1439460 $Y=1939440
X657 2 5217 5212 5252 3 NOR2X1 $T=1440780 1924720 1 0 $X=1440778 $Y=1919280
X658 2 5368 5342 5341 3 NOR2X1 $T=1459260 1934800 1 180 $X=1457280 $Y=1934398
X659 2 366 5339 5342 3 NOR2X1 $T=1459920 1965040 0 180 $X=1457940 $Y=1959600
X660 2 5445 5440 5426 3 NOR2X1 $T=1483020 1924720 1 180 $X=1481040 $Y=1924318
X661 2 379 384 5472 3 NOR2X1 $T=1486320 1985200 0 0 $X=1486318 $Y=1984798
X662 2 5474 5472 5501 3 NOR2X1 $T=1492920 1934800 0 0 $X=1492918 $Y=1934398
X663 2 391 389 5474 3 NOR2X1 $T=1494900 1965040 1 180 $X=1492920 $Y=1964638
X664 2 408 381 409 3 NOR2X1 $T=1519320 1783600 1 0 $X=1519318 $Y=1778160
X665 2 405 401 5612 3 NOR2X1 $T=1519320 1985200 1 0 $X=1519318 $Y=1979760
X666 2 358 363 5651 3 NOR2X1 $T=1521960 1793680 1 0 $X=1521958 $Y=1788240
X667 2 5609 5612 5561 3 NOR2X1 $T=1526580 1944880 1 180 $X=1524600 $Y=1944478
X668 2 410 407 5609 3 NOR2X1 $T=1527900 1965040 1 180 $X=1525920 $Y=1964638
X669 2 5746 414 5692 3 NOR2X1 $T=1532520 1934800 0 0 $X=1532518 $Y=1934398
X670 2 421 420 5715 3 NOR2X1 $T=1548360 1954960 0 0 $X=1548358 $Y=1954558
X671 2 5821 5805 5837 3 NOR2X1 $T=1556940 1884400 0 0 $X=1556938 $Y=1883998
X672 2 5864 5839 5838 3 NOR2X1 $T=1570800 1924720 1 180 $X=1568820 $Y=1924318
X673 2 5846 5802 5912 3 NOR2X1 $T=1582020 1894480 1 0 $X=1582018 $Y=1889040
X674 2 5883 443 5808 3 NOR2X1 $T=1591920 1783600 0 0 $X=1591918 $Y=1783198
X675 2 6326 478 6291 3 NOR2X1 $T=1682340 1904560 1 0 $X=1682338 $Y=1899120
X676 2 6442 491 6447 3 NOR2X1 $T=1699500 1954960 1 0 $X=1699498 $Y=1949520
X677 2 6518 497 6446 3 NOR2X1 $T=1718640 1924720 1 180 $X=1716660 $Y=1924318
X678 2 606 7235 7426 3 NOR2X1 $T=1917960 1965040 1 0 $X=1917958 $Y=1959600
X679 2 473 7609 7613 3 NOR2X1 $T=1976700 1823920 0 0 $X=1976698 $Y=1823518
X680 2 636 7683 7620 3 NOR2X1 $T=1997160 1884400 0 180 $X=1995180 $Y=1878960
X681 2 7782 7762 7744 3 NOR2X1 $T=2009040 1844080 1 180 $X=2007060 $Y=1843678
X682 2 7776 7783 7851 3 NOR2X1 $T=2029500 1985200 1 0 $X=2029498 $Y=1979760
X683 2 7840 7879 656 3 NOR2X1 $T=2042700 1965040 0 0 $X=2042698 $Y=1964638
X684 2 7851 656 7880 3 NOR2X1 $T=2044680 1985200 1 0 $X=2044678 $Y=1979760
X685 2 639 7837 7960 3 NOR2X1 $T=2048640 1823920 1 0 $X=2048638 $Y=1818480
X686 2 7547 663 7978 3 NOR2X1 $T=2065140 1783600 0 180 $X=2063160 $Y=1778160
X687 2 672 669 8054 3 NOR2X1 $T=2081640 1884400 0 180 $X=2079660 $Y=1878960
X688 2 7977 8001 670 3 NOR2X1 $T=2083620 1783600 1 0 $X=2083618 $Y=1778160
X689 2 7881 8039 8075 3 NOR2X1 $T=2085600 1975120 1 0 $X=2085598 $Y=1969680
X690 2 8052 8091 8107 3 NOR2X1 $T=2089560 1965040 1 0 $X=2089558 $Y=1959600
X691 2 8075 8107 8117 3 NOR2X1 $T=2092200 1985200 1 0 $X=2092198 $Y=1979760
X692 2 684 685 8182 3 NOR2X1 $T=2114640 1834000 1 0 $X=2114638 $Y=1828560
X693 2 8211 8273 693 3 NOR2X1 $T=2128500 1944880 1 0 $X=2128498 $Y=1939440
X694 2 8314 693 8307 3 NOR2X1 $T=2130480 1965040 1 180 $X=2128500 $Y=1964638
X695 2 8310 8288 8314 3 NOR2X1 $T=2140380 1965040 1 0 $X=2140378 $Y=1959600
X696 2 625 639 8308 3 NOR2X1 $T=2149620 1783600 0 0 $X=2149618 $Y=1783198
X697 2 8315 8365 711 3 NOR2X1 $T=2162820 1985200 0 0 $X=2162818 $Y=1984798
X698 2 8397 8495 8504 3 NOR2X1 $T=2189880 1954960 1 0 $X=2189878 $Y=1949520
X699 2 8496 708 8532 3 NOR2X1 $T=2195820 1834000 0 180 $X=2193840 $Y=1828560
X700 2 8512 8541 8596 3 NOR2X1 $T=2195160 1965040 0 0 $X=2195158 $Y=1964638
X701 2 711 8504 8624 3 NOR2X1 $T=2200440 1985200 1 0 $X=2200438 $Y=1979760
X702 2 8596 8600 8619 3 NOR2X1 $T=2205720 1975120 1 0 $X=2205718 $Y=1969680
X703 2 8582 8584 8600 3 NOR2X1 $T=2208360 1944880 1 180 $X=2206380 $Y=1944478
X704 2 8778 8869 8905 3 NOR2X1 $T=2276340 1884400 0 0 $X=2276338 $Y=1883998
X705 2 8889 8783 8996 3 NOR2X1 $T=2284260 1894480 0 0 $X=2284258 $Y=1894078
X706 2 8599 8798 8992 3 NOR2X1 $T=2289540 1944880 1 0 $X=2289538 $Y=1939440
X707 2 8800 8776 8983 3 NOR2X1 $T=2293500 1864240 1 0 $X=2293498 $Y=1858800
X708 2 8777 8814 9032 3 NOR2X1 $T=2304720 1944880 1 0 $X=2304718 $Y=1939440
X709 2 8983 8995 9024 3 NOR2X1 $T=2306700 1854160 0 0 $X=2306698 $Y=1853758
X710 2 8905 8996 9000 3 NOR2X1 $T=2306700 1884400 0 0 $X=2306698 $Y=1883998
X711 2 8797 8833 9068 3 NOR2X1 $T=2308680 1914640 1 0 $X=2308678 $Y=1909200
X712 2 8795 8832 9044 3 NOR2X1 $T=2311980 1924720 0 0 $X=2311978 $Y=1924318
X713 2 8992 9032 9113 3 NOR2X1 $T=2324520 1944880 1 0 $X=2324518 $Y=1939440
X714 2 9044 9068 9121 3 NOR2X1 $T=2327160 1924720 0 0 $X=2327158 $Y=1924318
X715 2 9163 9138 9191 3 NOR2X1 $T=2361480 1874320 1 0 $X=2361478 $Y=1868880
X716 2 9527 9454 9401 3 NOR2X1 $T=2401740 1944880 0 180 $X=2399760 $Y=1939440
X717 2 9475 9496 9517 3 NOR2X1 $T=2410980 1954960 1 0 $X=2410978 $Y=1949520
X718 2 9500 9497 9568 3 NOR2X1 $T=2420220 1834000 0 0 $X=2420218 $Y=1833598
X719 2 9707 9708 9761 3 NOR2X1 $T=2465760 1874320 1 0 $X=2465758 $Y=1868880
X720 2 792 799 9922 3 NOR2X1 $T=2490180 1985200 0 0 $X=2490178 $Y=1984798
X721 2 9836 9831 9921 3 NOR2X1 $T=2512620 1884400 0 180 $X=2510640 $Y=1878960
X722 2 10088 819 10065 3 NOR2X1 $T=2533740 1944880 0 180 $X=2531760 $Y=1939440
X723 2 826 827 10229 3 NOR2X1 $T=2544300 1793680 1 0 $X=2544298 $Y=1788240
X724 2 738 825 10119 3 NOR2X1 $T=2546280 1985200 1 180 $X=2544300 $Y=1984798
X725 2 10231 10233 10219 3 NOR2X1 $T=2562120 1914640 1 180 $X=2560140 $Y=1914238
X726 2 10248 830 10231 3 NOR2X1 $T=2562780 1944880 1 180 $X=2560800 $Y=1944478
X727 2 10252 10233 10217 3 NOR2X1 $T=2570700 1934800 1 0 $X=2570698 $Y=1929360
X728 2 828 10216 10300 3 NOR2X1 $T=2573340 1813840 1 0 $X=2573338 $Y=1808400
X729 2 834 832 10303 3 NOR2X1 $T=2579280 1975120 0 0 $X=2579278 $Y=1974718
X730 2 10229 10300 10339 3 NOR2X1 $T=2583900 1803760 0 0 $X=2583898 $Y=1803358
X731 59 1845 3 2 1814 NOR2X2 $T=688380 1793680 1 180 $X=685080 $Y=1793278
X732 1912 1963 3 2 65 NOR2X2 $T=711480 1793680 1 180 $X=708180 $Y=1793278
X733 65 1814 3 2 1974 NOR2X2 $T=711480 1793680 1 0 $X=711478 $Y=1788240
X734 1998 1975 3 2 2071 NOR2X2 $T=742500 1823920 1 0 $X=742498 $Y=1818480
X735 2063 2086 3 2 2070 NOR2X2 $T=748440 1944880 1 180 $X=745140 $Y=1944478
X736 2071 1997 3 2 73 NOR2X2 $T=750420 1803760 0 180 $X=747120 $Y=1798320
X737 75 77 3 2 2086 NOR2X2 $T=751740 1975120 1 180 $X=748440 $Y=1974718
X738 86 2195 3 2 2197 NOR2X2 $T=771540 1985200 0 180 $X=768240 $Y=1979760
X739 2363 2320 3 2 2297 NOR2X2 $T=799260 1803760 0 0 $X=799258 $Y=1803358
X740 2491 2469 3 2 2488 NOR2X2 $T=839520 1884400 0 180 $X=836220 $Y=1878960
X741 5168 4923 3 2 343 NOR2X2 $T=1422960 1834000 0 0 $X=1422958 $Y=1833598
X742 5439 5521 3 2 392 NOR2X2 $T=1494900 1783600 1 0 $X=1494898 $Y=1778160
X743 5795 5797 3 2 5687 NOR2X2 $T=1552980 1783600 1 180 $X=1549680 $Y=1783198
X744 424 5806 3 2 5795 NOR2X2 $T=1560240 1783600 0 0 $X=1560238 $Y=1783198
X745 468 6156 3 2 6119 NOR2X2 $T=1647360 1793680 1 0 $X=1647358 $Y=1788240
X746 7168 7167 3 2 6522 NOR2X2 $T=1868460 1834000 0 0 $X=1868458 $Y=1833598
X747 721 723 3 2 8625 NOR2X2 $T=2216940 1793680 1 0 $X=2216938 $Y=1788240
X748 742 8981 3 2 8979 NOR2X2 $T=2304060 1985200 0 180 $X=2300760 $Y=1979760
X749 9156 9142 3 2 754 NOR2X2 $T=2340360 1975120 0 180 $X=2337060 $Y=1969680
X750 10409 10412 3 2 10304 NOR2X2 $T=2601720 1793680 0 180 $X=2598420 $Y=1788240
X751 4612 4613 3 2 4610 OR2XL $T=1304160 1844080 1 180 $X=1301520 $Y=1843678
X752 417 418 3 2 411 OR2XL $T=1538460 1975120 0 180 $X=1535820 $Y=1969680
X753 6256 6251 3 2 6236 OR2XL $T=1662540 1944880 0 180 $X=1659900 $Y=1939440
X754 530 6787 3 2 6810 OR2XL $T=1790580 1793680 1 0 $X=1790578 $Y=1788240
X755 532 6863 3 2 6893 OR2XL $T=1803780 1844080 1 0 $X=1803778 $Y=1838640
X756 7439 7367 3 2 7566 OR2XL $T=1958220 1854160 0 0 $X=1958218 $Y=1853758
X757 532 713 3 2 8725 OR2XL $T=2232780 1874320 1 0 $X=2232778 $Y=1868880
X758 6753 725 3 2 8773 OR2XL $T=2238060 1854160 0 0 $X=2238058 $Y=1853758
X759 719 707 3 2 730 OR2XL $T=2240700 1783600 1 0 $X=2240698 $Y=1778160
X760 550 729 3 2 8816 OR2XL $T=2240700 1793680 1 0 $X=2240698 $Y=1788240
X761 557 725 3 2 8726 OR2XL $T=2244000 1894480 0 180 $X=2241360 $Y=1889040
X762 2034 2049 69 3 2 NAND2X2 $T=737880 1793680 1 180 $X=734580 $Y=1793278
X763 1974 73 2024 3 2 NAND2X2 $T=737880 1783600 0 0 $X=737878 $Y=1783198
X764 2917 2874 2894 3 2 NAND2X2 $T=931260 1803760 0 180 $X=927960 $Y=1798320
X765 3099 3137 3083 3 2 NAND2X2 $T=978120 1864240 1 180 $X=974820 $Y=1863838
X766 199 207 3715 3 2 NAND2X2 $T=1118700 1934800 1 0 $X=1118698 $Y=1929360
X767 4615 4500 4561 3 2 NAND2X2 $T=1296900 1813840 0 180 $X=1293600 $Y=1808400
X768 357 360 5216 3 2 NAND2X2 $T=1452000 1783600 1 180 $X=1448700 $Y=1783198
X769 369 360 5357 3 2 NAND2X2 $T=1465860 1783600 1 0 $X=1465858 $Y=1778160
X770 382 323 5453 3 2 NAND2X2 $T=1483020 1894480 1 0 $X=1483018 $Y=1889040
X771 402 5645 5671 3 2 NAND2X2 $T=1527240 1793680 1 0 $X=1527238 $Y=1788240
X772 5687 5685 5439 3 2 NAND2X2 $T=1531860 1783600 0 0 $X=1531858 $Y=1783198
X773 423 5806 5741 3 2 NAND2X2 $T=1553640 1783600 0 180 $X=1550340 $Y=1778160
X774 502 6559 6557 3 2 NAND2X2 $T=1732500 1844080 1 0 $X=1732498 $Y=1838640
X775 505 6576 6556 3 2 NAND2X2 $T=1738440 1854160 0 180 $X=1735140 $Y=1848720
X776 508 510 6544 3 2 NAND2X2 $T=1743060 1884400 1 0 $X=1743058 $Y=1878960
X777 6882 6803 6879 3 2 NAND2X2 $T=1807080 1975120 1 180 $X=1803780 $Y=1974718
X778 577 576 6926 3 2 NAND2X2 $T=1821600 1965040 1 180 $X=1818300 $Y=1964638
X779 583 7003 7004 3 2 NAND2X2 $T=1840080 1934800 1 180 $X=1836780 $Y=1934398
X780 600 599 602 3 2 NAND2X2 $T=1867140 1793680 1 0 $X=1867138 $Y=1788240
X781 605 7222 7204 3 2 NAND2X2 $T=1874400 1954960 1 180 $X=1871100 $Y=1954558
X782 8999 8976 749 3 2 NAND2X2 $T=2307360 1803760 1 0 $X=2307358 $Y=1798320
X783 9625 9459 9599 3 2 NAND2X2 $T=2442660 1914640 1 180 $X=2439360 $Y=1914238
X784 2154 2 2070 2137 3 2025 AOI21X4 $T=759000 1944880 0 180 $X=752400 $Y=1939440
X785 2471 2 2475 2465 3 2364 AOI21X4 $T=836220 1954960 0 180 $X=829620 $Y=1949520
X786 2916 2 2913 2902 3 2899 AOI21X4 $T=936540 1854160 1 180 $X=929940 $Y=1853758
X787 3789 2 46 4121 3 245 AOI21X4 $T=1203840 1783600 1 0 $X=1203838 $Y=1778160
X788 4615 2 4555 4629 3 4614 AOI21X4 $T=1302840 1813840 0 0 $X=1302838 $Y=1813438
X789 341 2 333 5203 3 347 AOI21X4 $T=1427580 1783600 1 0 $X=1427578 $Y=1778160
X790 7880 2 638 7883 3 7902 AOI21X4 $T=2034780 1985200 1 0 $X=2034778 $Y=1979760
X791 747 2 8976 8930 3 8937 AOI21X4 $T=2302080 1803760 0 180 $X=2295480 $Y=1798320
X792 8999 2 8930 9018 3 750 AOI21X4 $T=2306040 1793680 0 0 $X=2306038 $Y=1793278
X793 9401 2 9393 9378 3 8980 AOI21X4 $T=2396460 1934800 1 180 $X=2389860 $Y=1934398
X794 9786 2 9838 9921 3 10000 AOI21X4 $T=2497440 1874320 1 0 $X=2497438 $Y=1868880
X795 849 2 10056 10413 3 10410 AOI21X4 $T=2606340 1985200 0 180 $X=2599740 $Y=1979760
X796 88 2 90 3 2278 AND2X2 $T=780120 1783600 1 0 $X=780118 $Y=1778160
X797 2214 2 2272 3 2362 AND2X2 $T=794640 1934800 0 0 $X=794638 $Y=1934398
X798 2500 2 105 3 2405 AND2X2 $T=837540 1783600 1 180 $X=834900 $Y=1783198
X799 2732 2 2750 3 2694 AND2X2 $T=891000 1934800 0 180 $X=888360 $Y=1929360
X800 3061 2 3095 3 3099 AND2X2 $T=974820 1854160 0 0 $X=974818 $Y=1853758
X801 3621 2 3650 3 3651 AND2X2 $T=1100220 1854160 0 0 $X=1100218 $Y=1853758
X802 4365 2 3760 3 262 AND2X2 $T=1249380 1783600 0 0 $X=1249378 $Y=1783198
X803 4610 2 4632 3 4493 AND2X2 $T=1304160 1834000 1 180 $X=1301520 $Y=1833598
X804 323 2 321 3 4924 AND2X2 $T=1376100 1894480 0 180 $X=1373460 $Y=1889040
X805 5106 2 4998 3 5147 AND2X2 $T=1411740 1944880 0 0 $X=1411738 $Y=1944478
X806 5341 2 5228 3 5440 AND2X2 $T=1459920 1924720 0 0 $X=1459918 $Y=1924318
X807 382 2 387 3 5500 AND2X2 $T=1494240 1803760 0 0 $X=1494238 $Y=1803358
X808 5501 2 5561 3 5564 AND2X2 $T=1516680 1934800 1 180 $X=1514040 $Y=1934398
X809 5501 2 5589 3 5615 AND2X2 $T=1523940 1914640 1 0 $X=1523938 $Y=1909200
X810 426 2 5796 3 5797 AND2X2 $T=1556280 1793680 0 180 $X=1553640 $Y=1788240
X811 6142 2 448 3 6156 AND2X2 $T=1642080 1793680 1 0 $X=1642078 $Y=1788240
X812 6236 2 6169 3 477 AND2X2 $T=1662540 1954960 1 0 $X=1662538 $Y=1949520
X813 6396 2 492 3 6449 AND2X2 $T=1701480 1985200 0 0 $X=1701478 $Y=1984798
X814 511 2 6599 3 506 AND2X2 $T=1740420 1954960 1 180 $X=1737780 $Y=1954558
X815 544 2 6813 3 6576 AND2X2 $T=1789260 1844080 1 180 $X=1786620 $Y=1843678
X816 526 2 7147 3 7168 AND2X2 $T=1862520 1834000 0 0 $X=1862518 $Y=1833598
X817 597 2 7234 3 7211 AND2X2 $T=1895520 1864240 1 180 $X=1892880 $Y=1863838
X818 7783 2 7776 3 7779 AND2X2 $T=2015640 1975120 1 180 $X=2013000 $Y=1974718
X819 639 2 625 3 8272 AND2X2 $T=2143680 1783600 1 0 $X=2143678 $Y=1778160
X820 8976 2 8904 3 8991 AND2X2 $T=2311320 1823920 0 180 $X=2308680 $Y=1818480
X821 9000 2 9024 3 9027 AND2X2 $T=2319240 1874320 1 180 $X=2316600 $Y=1873918
X822 9026 2 9129 3 9084 AND2X2 $T=2337720 1874320 1 180 $X=2335080 $Y=1873918
X823 9540 2 9456 3 9496 AND2X2 $T=2420880 1954960 0 180 $X=2418240 $Y=1949520
X824 9707 2 9708 3 9775 AND2X2 $T=2464440 1864240 1 0 $X=2464438 $Y=1858800
X825 807 2 9922 3 9973 AND2X2 $T=2515260 1985200 0 0 $X=2515258 $Y=1984798
X826 3063 3 3083 2 2916 NAND2X4 $T=972180 1864240 1 180 $X=967560 $Y=1863838
X827 5466 3 322 2 380 NAND2X4 $T=1484340 1884400 0 180 $X=1479720 $Y=1878960
X828 5570 3 5585 2 357 NAND2X4 $T=1504140 1793680 1 0 $X=1504138 $Y=1788240
X829 447 3 5973 2 446 NAND2X4 $T=1599840 1864240 0 180 $X=1595220 $Y=1858800
X830 148 3 457 2 6066 NAND2X4 $T=1618980 1793680 0 0 $X=1618978 $Y=1793278
X831 2071 2050 3 2 2034 OR2X2 $T=739860 1803760 1 180 $X=737220 $Y=1803358
X832 2291 2275 3 2 2214 OR2X2 $T=792000 1965040 0 180 $X=789360 $Y=1959600
X833 2297 2294 3 2 92 OR2X2 $T=793320 1823920 1 180 $X=790680 $Y=1823518
X834 2732 2750 3 2 2699 OR2X2 $T=894960 1944880 0 180 $X=892320 $Y=1939440
X835 2315 120 3 2 2913 OR2X2 $T=937200 1854160 0 180 $X=934560 $Y=1848720
X836 50 62 3 2 2935 OR2X2 $T=937200 1934800 0 0 $X=937198 $Y=1934398
X837 2841 3212 3 2 3095 OR2X2 $T=1005180 1864240 1 180 $X=1002540 $Y=1863838
X838 2842 3321 3 2 3298 OR2X2 $T=1034880 1904560 1 0 $X=1034878 $Y=1899120
X839 176 177 3 2 3463 OR2X2 $T=1073160 1813840 0 0 $X=1073158 $Y=1813438
X840 3514 3513 3 2 3526 OR2X2 $T=1084380 1904560 0 180 $X=1081740 $Y=1899120
X841 179 187 3 2 3522 OR2X2 $T=1084380 1975120 0 0 $X=1084378 $Y=1974718
X842 196 168 3 2 195 OR2X2 $T=1089660 1985200 1 180 $X=1087020 $Y=1984798
X843 198 199 3 2 3621 OR2X2 $T=1097580 1854160 1 0 $X=1097578 $Y=1848720
X844 3622 3651 3 2 3657 OR2X2 $T=1100220 1874320 0 0 $X=1100218 $Y=1873918
X845 204 205 3 2 3654 OR2X2 $T=1117380 1823920 1 180 $X=1114740 $Y=1823518
X846 3453 206 3 2 3738 OR2X2 $T=1117380 1854160 0 0 $X=1117378 $Y=1853758
X847 3918 3931 3 2 3880 OR2X2 $T=1166880 1844080 0 180 $X=1164240 $Y=1838640
X848 4033 4025 3 2 3970 OR2X2 $T=1189320 1884400 0 180 $X=1186680 $Y=1878960
X849 3431 4117 3 2 4127 OR2X2 $T=1201200 1914640 0 0 $X=1201198 $Y=1914238
X850 4128 4124 3 2 4047 OR2X2 $T=1205160 1864240 1 180 $X=1202520 $Y=1863838
X851 4312 4288 3 2 4256 OR2X2 $T=1236180 1874320 0 180 $X=1233540 $Y=1868880
X852 3589 4327 3 2 4314 OR2X2 $T=1244100 1914640 1 180 $X=1241460 $Y=1914238
X853 4453 4489 3 2 4433 OR2X2 $T=1278420 1884400 0 180 $X=1275780 $Y=1878960
X854 3010 4495 3 2 4500 OR2X2 $T=1278420 1834000 1 0 $X=1278418 $Y=1828560
X855 266 68 3 2 4474 OR2X2 $T=1281060 1834000 1 180 $X=1278420 $Y=1833598
X856 3832 4503 3 2 4483 OR2X2 $T=1282380 1904560 1 180 $X=1279740 $Y=1904158
X857 4485 286 3 2 4609 OR2X2 $T=1300200 1874320 1 0 $X=1300198 $Y=1868880
X858 4918 4921 3 2 4929 OR2X2 $T=1372140 1854160 1 0 $X=1372138 $Y=1848720
X859 4923 5028 3 2 5083 OR2X2 $T=1398540 1834000 0 0 $X=1398538 $Y=1833598
X860 368 374 3 2 5403 OR2X2 $T=1473120 1975120 0 0 $X=1473118 $Y=1974718
X861 398 399 3 2 5586 OR2X2 $T=1504140 1844080 0 0 $X=1504138 $Y=1843678
X862 5765 5772 3 2 5798 OR2X2 $T=1550340 1934800 1 0 $X=1550338 $Y=1929360
X863 5837 5838 3 2 5846 OR2X2 $T=1563540 1884400 0 0 $X=1563538 $Y=1883998
X864 5939 5951 3 2 5935 OR2X2 $T=1594560 1904560 0 180 $X=1591920 $Y=1899120
X865 5932 5921 3 2 5974 OR2X2 $T=1602480 1924720 1 0 $X=1602478 $Y=1919280
X866 464 6083 3 2 6080 OR2X2 $T=1626240 1975120 1 180 $X=1623600 $Y=1974718
X867 473 111 3 2 6249 OR2X2 $T=1659900 1844080 1 0 $X=1659898 $Y=1838640
X868 479 6333 3 2 6296 OR2X2 $T=1683660 1965040 0 0 $X=1683658 $Y=1964638
X869 486 6377 3 2 6294 OR2X2 $T=1699500 1924720 1 0 $X=1699498 $Y=1919280
X870 494 6451 3 2 6464 OR2X2 $T=1703460 1975120 0 0 $X=1703458 $Y=1974718
X871 516 517 3 2 6678 OR2X2 $T=1756920 1944880 0 0 $X=1756918 $Y=1944478
X872 6678 319 3 2 525 OR2X2 $T=1767480 1934800 1 0 $X=1767478 $Y=1929360
X873 6678 310 3 2 556 OR2X2 $T=1773420 1965040 1 0 $X=1773418 $Y=1959600
X874 6678 303 3 2 540 OR2X2 $T=1780680 1934800 1 0 $X=1780678 $Y=1929360
X875 6678 308 3 2 543 OR2X2 $T=1780680 1944880 1 0 $X=1780678 $Y=1939440
X876 6660 549 3 2 548 OR2X2 $T=1797180 1954960 0 180 $X=1794540 $Y=1949520
X877 6660 551 3 2 555 OR2X2 $T=1797180 1944880 1 0 $X=1797178 $Y=1939440
X878 553 558 3 2 6803 OR2X2 $T=1803780 1975120 1 0 $X=1803778 $Y=1969680
X879 6660 566 3 2 563 OR2X2 $T=1813020 1944880 0 180 $X=1810380 $Y=1939440
X880 6660 567 3 2 569 OR2X2 $T=1811700 1954960 1 0 $X=1811698 $Y=1949520
X881 7468 622 3 2 7406 OR2X2 $T=1950300 1894480 1 180 $X=1947660 $Y=1894078
X882 7407 611 3 2 7470 OR2X2 $T=1958220 1944880 1 180 $X=1955580 $Y=1944478
X883 7543 625 3 2 7527 OR2X2 $T=1963500 1934800 1 180 $X=1960860 $Y=1934398
X884 7591 7234 3 2 7616 OR2X2 $T=1978020 1954960 1 0 $X=1978018 $Y=1949520
X885 7657 629 3 2 7573 OR2X2 $T=1983300 1904560 0 180 $X=1980660 $Y=1899120
X886 7699 7679 3 2 7643 OR2X2 $T=1995840 1954960 1 180 $X=1993200 $Y=1954558
X887 648 644 3 2 7800 OR2X2 $T=2028840 1874320 0 180 $X=2026200 $Y=1868880
X888 642 625 3 2 7852 OR2X2 $T=2028840 1783600 1 0 $X=2028838 $Y=1778160
X889 654 653 3 2 7861 OR2X2 $T=2042700 1894480 0 180 $X=2040060 $Y=1889040
X890 681 680 3 2 8119 OR2X2 $T=2103420 1864240 0 180 $X=2100780 $Y=1858800
X891 8212 8096 3 2 8189 OR2X2 $T=2112660 1944880 1 180 $X=2110020 $Y=1944478
X892 8921 8920 3 2 741 OR2X2 $T=2292840 1985200 0 180 $X=2290200 $Y=1979760
X893 8779 8831 3 2 9031 OR2X2 $T=2298120 1834000 1 0 $X=2298118 $Y=1828560
X894 8780 8939 3 2 9023 OR2X2 $T=2298120 1844080 0 0 $X=2298118 $Y=1843678
X895 8812 9042 3 2 748 OR2X2 $T=2316600 1975120 0 180 $X=2313960 $Y=1969680
X896 9120 9137 3 2 8976 OR2X2 $T=2341680 1823920 0 180 $X=2339040 $Y=1818480
X897 9269 9241 3 2 9242 OR2X2 $T=2367420 1965040 0 0 $X=2367418 $Y=1964638
X898 9114 9302 3 2 9317 OR2X2 $T=2374020 1934800 1 0 $X=2374018 $Y=1929360
X899 9318 9316 3 2 9346 OR2X2 $T=2395140 1965040 0 180 $X=2392500 $Y=1959600
X900 9472 9458 3 2 9457 OR2X2 $T=2406360 1874320 1 180 $X=2403720 $Y=1873918
X901 9625 9459 3 2 9627 OR2X2 $T=2440680 1924720 0 0 $X=2440678 $Y=1924318
X902 9759 9811 3 2 9794 OR2X2 $T=2488200 1844080 1 0 $X=2488198 $Y=1838640
X903 10231 10065 3 2 10252 OR2X2 $T=2564760 1944880 1 0 $X=2564758 $Y=1939440
X904 10254 10231 3 2 10268 OR2X2 $T=2583240 1914640 1 180 $X=2580600 $Y=1914238
X905 30 3 2 27 19 NAND2XL $T=663300 1985200 0 180 $X=661320 $Y=1979760
X906 24 3 2 42 1757 NAND2XL $T=671220 1924720 1 180 $X=669240 $Y=1924318
X907 3045 3 2 3061 3098 NAND2XL $T=972840 1854160 1 0 $X=972838 $Y=1848720
X908 3324 3 2 3298 3358 NAND2XL $T=1035540 1914640 0 0 $X=1035538 $Y=1914238
X909 177 3 2 176 3452 NAND2XL $T=1065900 1823920 1 180 $X=1063920 $Y=1823518
X910 3674 3 2 3654 3615 NAND2XL $T=1105500 1823920 1 180 $X=1103520 $Y=1823518
X911 206 3 2 3453 3734 NAND2XL $T=1117380 1864240 0 0 $X=1117378 $Y=1863838
X912 3734 3 2 3738 3814 NAND2XL $T=1131240 1864240 1 0 $X=1131238 $Y=1858800
X913 3913 3 2 3880 3811 NAND2XL $T=1155000 1834000 0 180 $X=1153020 $Y=1828560
X914 4013 3 2 3970 3969 NAND2XL $T=1184040 1864240 0 180 $X=1182060 $Y=1858800
X915 4030 3 2 3475 4003 NAND2XL $T=1188000 1914640 0 0 $X=1187998 $Y=1914238
X916 4178 3 2 4126 4079 NAND2XL $T=1205820 1874320 1 180 $X=1203840 $Y=1873918
X917 4231 3 2 4199 4240 NAND2XL $T=1224960 1944880 1 0 $X=1224958 $Y=1939440
X918 4287 3 2 4256 4260 NAND2XL $T=1233540 1854160 1 180 $X=1231560 $Y=1853758
X919 4304 3 2 4314 4348 NAND2XL $T=1242120 1914640 1 0 $X=1242118 $Y=1909200
X920 4417 3 2 4433 4439 NAND2XL $T=1262580 1884400 1 0 $X=1262578 $Y=1878960
X921 68 3 2 266 3897 NAND2XL $T=1265220 1844080 1 0 $X=1265218 $Y=1838640
X922 4501 3 2 4500 4471 NAND2XL $T=1280400 1813840 1 180 $X=1278420 $Y=1813438
X923 4533 3 2 4483 4539 NAND2XL $T=1287660 1904560 1 0 $X=1287658 $Y=1899120
X924 4550 3 2 4532 4516 NAND2XL $T=1295580 1884400 0 180 $X=1293600 $Y=1878960
X925 4684 3 2 3933 4673 NAND2XL $T=1322640 1894480 0 180 $X=1320660 $Y=1889040
X926 4615 3 2 4693 4687 NAND2XL $T=1325940 1813840 1 0 $X=1325938 $Y=1808400
X927 4746 3 2 4706 4765 NAND2XL $T=1338480 1834000 1 0 $X=1338478 $Y=1828560
X928 4930 3 2 4915 4949 NAND2XL $T=1375440 1944880 1 0 $X=1375438 $Y=1939440
X929 328 3 2 327 4967 NAND2XL $T=1391940 1965040 1 180 $X=1389960 $Y=1964638
X930 5104 3 2 5027 5080 NAND2XL $T=1400520 1854160 0 180 $X=1398540 $Y=1848720
X931 5199 3 2 5236 5202 NAND2XL $T=1441440 1954960 0 180 $X=1439460 $Y=1949520
X932 5252 3 2 5324 5343 NAND2XL $T=1453980 1914640 0 0 $X=1453978 $Y=1914238
X933 5442 3 2 5467 5425 NAND2XL $T=1481700 1904560 1 180 $X=1479720 $Y=1904158
X934 391 3 2 389 5438 NAND2XL $T=1496220 1975120 0 180 $X=1494240 $Y=1969680
X935 5581 3 2 5589 5563 NAND2XL $T=1505460 1914640 0 180 $X=1503480 $Y=1909200
X936 5501 3 2 5523 5588 NAND2XL $T=1513380 1914640 0 180 $X=1511400 $Y=1909200
X937 5615 3 2 5523 5633 NAND2XL $T=1523940 1904560 1 180 $X=1521960 $Y=1904158
X938 5821 3 2 5805 5841 NAND2XL $T=1556940 1894480 1 0 $X=1556938 $Y=1889040
X939 5864 3 2 5839 5862 NAND2XL $T=1573440 1924720 1 180 $X=1571460 $Y=1924318
X940 6083 3 2 464 6129 NAND2XL $T=1636800 1975120 0 0 $X=1636798 $Y=1974718
X941 111 3 2 473 474 NAND2XL $T=1660560 1823920 0 0 $X=1660558 $Y=1823518
X942 6326 3 2 478 6276 NAND2XL $T=1672440 1904560 0 180 $X=1670460 $Y=1899120
X943 6293 3 2 6296 6315 NAND2XL $T=1673760 1965040 1 0 $X=1673758 $Y=1959600
X944 6442 3 2 491 6450 NAND2XL $T=1702140 1954960 1 0 $X=1702138 $Y=1949520
X945 6501 3 2 6464 6502 NAND2XL $T=1719960 1975120 1 180 $X=1717980 $Y=1974718
X946 6518 3 2 497 6448 NAND2XL $T=1721280 1934800 1 180 $X=1719300 $Y=1934398
X947 6812 3 2 6803 546 NAND2XL $T=1793220 1985200 0 180 $X=1791240 $Y=1979760
X948 6926 3 2 6882 6782 NAND2XL $T=1828200 1975120 0 180 $X=1826220 $Y=1969680
X949 559 3 2 7367 7350 NAND2XL $T=1928520 1844080 0 0 $X=1928518 $Y=1843678
X950 7403 3 2 7406 7417 NAND2XL $T=1934460 1894480 0 0 $X=1934458 $Y=1894078
X951 622 3 2 7468 7403 NAND2XL $T=1945020 1894480 1 180 $X=1943040 $Y=1894078
X952 7472 3 2 7470 7440 NAND2XL $T=1948980 1954960 1 180 $X=1947000 $Y=1954558
X953 7525 3 2 7527 7422 NAND2XL $T=1958220 1975120 1 180 $X=1956240 $Y=1974718
X954 7646 3 2 7573 7526 NAND2XL $T=1978680 1894480 1 180 $X=1976700 $Y=1894078
X955 7660 3 2 7643 7644 NAND2XL $T=1986600 1965040 0 180 $X=1984620 $Y=1959600
X956 7799 3 2 7800 7637 NAND2XL $T=2011680 1874320 0 180 $X=2009700 $Y=1868880
X957 7818 3 2 7817 7821 NAND2XL $T=2034120 1803760 1 180 $X=2032140 $Y=1803358
X958 625 3 2 642 7929 NAND2XL $T=2049960 1783600 1 0 $X=2049958 $Y=1778160
X959 8006 3 2 7976 7921 NAND2XL $T=2058540 1864240 1 180 $X=2056560 $Y=1863838
X960 659 3 2 661 8006 NAND2XL $T=2065140 1864240 1 0 $X=2065138 $Y=1858800
X961 8169 3 2 8119 8057 NAND2XL $T=2093520 1864240 0 180 $X=2091540 $Y=1858800
X962 8233 3 2 8189 8190 NAND2XL $T=2117940 1975120 1 0 $X=2117938 $Y=1969680
X963 721 3 2 723 8612 NAND2XL $T=2211660 1793680 0 180 $X=2209680 $Y=1788240
X964 8778 3 2 8869 8919 NAND2XL $T=2276340 1874320 0 0 $X=2276338 $Y=1873918
X965 9052 3 2 8999 8982 NAND2XL $T=2319900 1803760 0 180 $X=2317920 $Y=1798320
X966 9072 3 2 9219 9220 NAND2XL $T=2350920 1934800 1 0 $X=2350918 $Y=1929360
X967 9245 3 2 9242 762 NAND2XL $T=2360820 1975120 1 180 $X=2358840 $Y=1974718
X968 8993 3 2 9240 9272 NAND2XL $T=2366760 1854160 0 0 $X=2366758 $Y=1853758
X969 9219 3 2 9113 9302 NAND2XL $T=2366760 1934800 1 0 $X=2366758 $Y=1929360
X970 9320 3 2 9346 769 NAND2XL $T=2384580 1975120 1 180 $X=2382600 $Y=1974718
X971 9473 3 2 9457 9453 NAND2XL $T=2402400 1914640 1 180 $X=2400420 $Y=1914238
X972 9455 3 2 9456 777 NAND2XL $T=2405700 1965040 1 0 $X=2405698 $Y=1959600
X973 9504 3 2 9494 9377 NAND2XL $T=2411640 1854160 1 180 $X=2409660 $Y=1853758
X974 9550 3 2 9593 9573 NAND2XL $T=2430120 1934800 0 180 $X=2428140 $Y=1929360
X975 9814 3 2 9794 9779 NAND2XL $T=2475660 1854160 1 180 $X=2473680 $Y=1853758
X976 9786 3 2 9838 9865 NAND2XL $T=2489520 1874320 1 0 $X=2489518 $Y=1868880
X977 839 3 2 840 845 NAND2XL $T=2583900 1783600 0 0 $X=2583898 $Y=1783198
X978 3434 3438 3 2 INVX4 $T=1058640 1965040 1 0 $X=1058638 $Y=1959600
X979 190 196 3 2 INVX4 $T=1092960 1944880 0 0 $X=1092958 $Y=1944478
X980 150 108 3 2 INVX4 $T=1111440 1793680 0 0 $X=1111438 $Y=1793278
X981 180 187 3 2 INVX4 $T=1120680 1975120 1 180 $X=1118040 $Y=1974718
X982 111 152 3 2 INVX4 $T=1134540 1813840 0 0 $X=1134538 $Y=1813438
X983 511 6695 3 2 INVX4 $T=1760220 1965040 1 0 $X=1760218 $Y=1959600
X984 7043 6983 3 2 INVX4 $T=1855920 1894480 0 0 $X=1855918 $Y=1894078
X985 521 7098 3 2 INVX4 $T=2101440 1894480 0 0 $X=2101438 $Y=1894078
X986 9393 9505 3 2 INVX4 $T=2413620 1975120 0 0 $X=2413618 $Y=1974718
X987 10082 10302 3 2 INVX4 $T=2586540 1823920 1 0 $X=2586538 $Y=1818480
X988 85 2195 2 2197 2208 3 AOI21X1 $T=774180 1975120 1 180 $X=771540 $Y=1974718
X989 2214 2279 2 2274 2271 3 AOI21X1 $T=789360 1934800 0 180 $X=786720 $Y=1929360
X990 2450 2447 2 2446 102 3 AOI21X1 $T=828300 1823920 0 180 $X=825660 $Y=1818480
X991 2693 2633 2 2588 2619 3 AOI21X1 $T=866580 1894480 0 180 $X=863940 $Y=1889040
X992 2699 2695 2 2694 2634 3 AOI21X1 $T=883080 1944880 0 180 $X=880440 $Y=1939440
X993 2664 2697 2 2693 2656 3 AOI21X1 $T=883740 1894480 1 180 $X=881100 $Y=1894078
X994 2749 2730 2 2727 2663 3 AOI21X1 $T=891000 1844080 0 180 $X=888360 $Y=1838640
X995 2935 2933 2 2930 2859 3 AOI21X1 $T=940500 1924720 1 180 $X=937860 $Y=1924318
X996 3061 3067 2 3062 3063 3 AOI21X1 $T=970200 1854160 1 180 $X=967560 $Y=1853758
X997 3121 3069 2 3064 2660 3 AOI21X1 $T=970200 1894480 0 180 $X=967560 $Y=1889040
X998 3095 3137 2 3067 3132 3 AOI21X1 $T=989340 1864240 0 180 $X=986700 $Y=1858800
X999 3322 3298 2 3295 3292 3 AOI21X1 $T=1030260 1904560 1 180 $X=1027620 $Y=1904158
X1000 182 3479 2 178 156 3 AOI21X1 $T=1071840 1783600 0 180 $X=1069200 $Y=1778160
X1001 3526 3495 2 3484 3366 3 AOI21X1 $T=1071840 1904560 1 180 $X=1069200 $Y=1904158
X1002 179 187 2 3504 3476 3 AOI21X1 $T=1077120 1975120 1 180 $X=1074480 $Y=1974718
X1003 3654 3610 2 3609 3567 3 AOI21X1 $T=1098900 1823920 1 180 $X=1096260 $Y=1823518
X1004 3735 3657 2 3698 3673 3 AOI21X1 $T=1118040 1894480 0 180 $X=1115400 $Y=1889040
X1005 3970 3972 2 3985 3807 3 AOI21X1 $T=1174140 1864240 0 0 $X=1174138 $Y=1863838
X1006 4127 4125 2 4122 4045 3 AOI21X1 $T=1205160 1914640 0 180 $X=1202520 $Y=1909200
X1007 4261 4256 2 4251 4124 3 AOI21X1 $T=1229580 1864240 0 180 $X=1226940 $Y=1858800
X1008 4314 4313 2 4310 4224 3 AOI21X1 $T=1242780 1904560 0 180 $X=1240140 $Y=1899120
X1009 4440 4433 2 4432 4366 3 AOI21X1 $T=1263900 1864240 1 180 $X=1261260 $Y=1863838
X1010 4486 4483 2 4480 4408 3 AOI21X1 $T=1277100 1904560 0 180 $X=1274460 $Y=1899120
X1011 4500 4470 2 4555 4635 3 AOI21X1 $T=1294920 1823920 1 0 $X=1294918 $Y=1818480
X1012 4915 4902 2 4901 4900 3 AOI21X1 $T=1368180 1944880 0 180 $X=1365540 $Y=1939440
X1013 4998 4902 2 4999 5009 3 AOI21X1 $T=1391940 1934800 1 0 $X=1391938 $Y=1929360
X1014 4999 5106 2 5108 5131 3 AOI21X1 $T=1407780 1944880 1 0 $X=1407778 $Y=1939440
X1015 5274 338 2 357 359 3 AOI21X1 $T=1448700 1793680 1 0 $X=1448698 $Y=1788240
X1016 6304 6296 2 6321 6349 3 AOI21X1 $T=1678380 1965040 1 0 $X=1678378 $Y=1959600
X1017 6292 6294 2 6361 6399 3 AOI21X1 $T=1687620 1924720 0 0 $X=1687618 $Y=1924318
X1018 6464 6482 2 6540 499 3 AOI21X1 $T=1725240 1975120 0 0 $X=1725238 $Y=1974718
X1019 521 527 2 545 6699 3 AOI21X1 $T=1791900 1834000 1 180 $X=1789260 $Y=1833598
X1020 6803 552 2 6821 6783 3 AOI21X1 $T=1797180 1985200 1 0 $X=1797178 $Y=1979760
X1021 6821 6882 2 6936 6899 3 AOI21X1 $T=1820280 1985200 1 0 $X=1820278 $Y=1979760
X1022 607 596 2 7211 7099 3 AOI21X1 $T=1882320 1864240 1 180 $X=1879680 $Y=1863838
X1023 7527 7421 2 7542 627 3 AOI21X1 $T=1960860 1975120 0 0 $X=1960858 $Y=1974718
X1024 7445 7573 2 7587 7586 3 AOI21X1 $T=1970100 1894480 0 0 $X=1970098 $Y=1894078
X1025 7616 7610 2 7619 7623 3 AOI21X1 $T=1979340 1965040 1 0 $X=1979338 $Y=1959600
X1026 7619 7643 2 7662 7684 3 AOI21X1 $T=1992540 1965040 1 0 $X=1992538 $Y=1959600
X1027 7800 7636 2 7813 7819 3 AOI21X1 $T=2020920 1874320 1 0 $X=2020918 $Y=1868880
X1028 7761 7817 2 7820 652 3 AOI21X1 $T=2023560 1803760 1 0 $X=2023558 $Y=1798320
X1029 8117 665 2 8130 8183 3 AOI21X1 $T=2096820 1985200 0 0 $X=2096818 $Y=1984798
X1030 8130 8189 2 8217 8218 3 AOI21X1 $T=2112660 1975120 1 0 $X=2112658 $Y=1969680
X1031 8602 8619 2 8623 8640 3 AOI21X1 $T=2211660 1975120 1 0 $X=2211658 $Y=1969680
X1032 8712 726 2 8717 8716 3 AOI21X1 $T=2238060 1975120 0 0 $X=2238058 $Y=1974718
X1033 9021 9024 2 9025 9039 3 AOI21X1 $T=2311320 1864240 1 0 $X=2311318 $Y=1858800
X1034 9129 9073 2 9075 9076 3 AOI21X1 $T=2327160 1874320 0 180 $X=2324520 $Y=1868880
X1035 9040 9121 2 9112 9116 3 AOI21X1 $T=2335080 1924720 0 180 $X=2332440 $Y=1919280
X1036 9109 9073 2 9157 9164 3 AOI21X1 $T=2340360 1894480 0 0 $X=2340358 $Y=1894078
X1037 9191 9073 2 9168 9174 3 AOI21X1 $T=2348280 1874320 0 180 $X=2345640 $Y=1868880
X1038 9113 8659 2 9040 9237 3 AOI21X1 $T=2355540 1934800 0 0 $X=2355538 $Y=1934398
X1039 9242 766 2 9287 767 3 AOI21X1 $T=2370060 1985200 1 0 $X=2370058 $Y=1979760
X1040 9346 9287 2 9371 9366 3 AOI21X1 $T=2387220 1975120 0 0 $X=2387218 $Y=1974718
X1041 9475 9457 2 9479 9483 3 AOI21X1 $T=2405700 1934800 1 0 $X=2405698 $Y=1929360
X1042 9762 9615 2 9775 9780 3 AOI21X1 $T=2469720 1874320 0 0 $X=2469718 $Y=1873918
X1043 9775 9794 2 9835 9838 3 AOI21X1 $T=2488200 1864240 1 0 $X=2488198 $Y=1858800
X1044 807 803 2 809 9974 3 AOI21X1 $T=2508660 1985200 0 0 $X=2508658 $Y=1984798
X1045 10056 10217 2 10215 10095 3 AOI21X1 $T=2554860 1934800 0 180 $X=2552220 $Y=1929360
X1046 10286 10056 2 10290 10255 3 AOI21X1 $T=2573340 1914640 1 0 $X=2573338 $Y=1909200
X1047 2136 2063 3 2051 2 2137 OAI21X2 $T=755040 1954960 0 180 $X=749760 $Y=1949520
X1048 92 2280 3 2250 2 94 OAI21X2 $T=789360 1813840 0 180 $X=784080 $Y=1808400
X1049 2299 2297 3 2361 2 82 OAI21X2 $T=796620 1823920 0 0 $X=796618 $Y=1823518
X1050 2480 2529 3 2451 2 2454 OAI21X2 $T=836880 1934800 1 180 $X=831600 $Y=1934398
X1051 3873 3807 3 3820 2 3810 OAI21X2 $T=1153020 1864240 0 0 $X=1153018 $Y=1863838
X1052 7698 7639 3 7684 2 638 OAI21X2 $T=2000460 1975120 0 180 $X=1995180 $Y=1969680
X1053 8089 8038 3 8129 2 8205 OAI21X2 $T=2094840 1803760 1 0 $X=2094838 $Y=1798320
X1054 8205 690 3 8281 2 8364 OAI21X2 $T=2127180 1813840 1 0 $X=2127178 $Y=1808400
X1055 8364 8393 3 8429 2 8444 OAI21X2 $T=2170080 1813840 1 180 $X=2164800 $Y=1813438
X1056 754 752 3 9094 2 756 OAI21X2 $T=2335740 1985200 1 0 $X=2335738 $Y=1979760
X1057 9594 9505 3 9599 2 9570 OAI21X2 $T=2431440 1975120 0 0 $X=2431438 $Y=1974718
X1058 10302 10300 3 10269 2 10270 OAI21X2 $T=2577960 1813840 0 0 $X=2577958 $Y=1813438
X1059 8991 8980 743 3 2 XNOR2X4 $T=2306700 1924720 0 180 $X=2295480 $Y=1919280
X1060 9726 791 794 3 2 XNOR2X4 $T=2458500 1965040 1 0 $X=2458498 $Y=1959600
X1061 815 10009 811 3 2 XNOR2X4 $T=2523840 1924720 1 180 $X=2512620 $Y=1924318
X1062 10360 10056 831 3 2 XNOR2X4 $T=2596440 1904560 1 180 $X=2585220 $Y=1904158
X1063 2025 3 2024 1993 2 70 OAI21X4 $T=733920 1783600 1 180 $X=726660 $Y=1783198
X1064 2364 3 2213 2205 2 2154 OAI21X4 $T=775500 1944880 1 180 $X=768240 $Y=1944478
X1065 2660 3 2638 2619 2 95 OAI21X4 $T=869880 1894480 1 180 $X=862620 $Y=1894078
X1066 2894 3 2899 2910 2 119 OAI21X4 $T=927960 1793680 1 0 $X=927958 $Y=1788240
X1067 4311 3 3962 4286 2 258 OAI21X4 $T=1241460 1823920 1 0 $X=1241458 $Y=1818480
X1068 4561 3 3991 4614 2 288 OAI21X4 $T=1300200 1803760 0 0 $X=1300198 $Y=1803358
X1069 5271 3 341 4863 2 5082 OAI21X4 $T=1417020 1783600 1 180 $X=1409760 $Y=1783198
X1070 6879 3 564 6899 2 571 OAI21X4 $T=1809720 1975120 0 0 $X=1809718 $Y=1974718
X1071 8054 3 8004 8056 2 8051 OAI21X4 $T=2076360 1874320 0 0 $X=2076358 $Y=1873918
X1072 8182 3 8115 8170 2 683 OAI21X4 $T=2106720 1834000 1 180 $X=2099460 $Y=1833598
X1073 8317 3 8660 8640 2 8659 OAI21X4 $T=2224200 1975120 0 180 $X=2216940 $Y=1969680
X1074 9321 3 770 9366 2 9393 OAI21X4 $T=2382600 1985200 0 0 $X=2382598 $Y=1984798
X1075 144 3 50 2 CLKBUFX8 $T=993300 1793680 1 0 $X=993298 $Y=1788240
X1076 4155 3 190 2 CLKBUFX8 $T=1212420 1954960 0 180 $X=1207800 $Y=1949520
X1077 300 3 68 2 CLKBUFX8 $T=1331220 1783600 1 180 $X=1326600 $Y=1783198
X1078 4880 3 230 2 CLKBUFX8 $T=1364880 1914640 0 180 $X=1360260 $Y=1909200
X1079 382 3 395 2 CLKBUFX8 $T=1492920 1864240 0 0 $X=1492918 $Y=1863838
X1080 7368 3 616 2 CLKBUFX8 $T=1923900 1793680 0 180 $X=1919280 $Y=1788240
X1081 624 3 623 2 CLKBUFX8 $T=1960860 1985200 1 180 $X=1956240 $Y=1984798
X1082 7569 3 625 2 CLKBUFX8 $T=1970760 1813840 0 180 $X=1966140 $Y=1808400
X1083 10214 3 829 2 CLKBUFX8 $T=2554200 1864240 1 180 $X=2549580 $Y=1863838
X1084 2134 2135 2 3 80 XOR2X2 $T=749760 1793680 1 0 $X=749758 $Y=1788240
X1085 2282 2280 2 3 2315 XOR2X2 $T=790020 1834000 0 0 $X=790018 $Y=1833598
X1086 2448 2454 2 3 2469 XOR2X2 $T=826980 1924720 0 0 $X=826978 $Y=1924318
X1087 7819 7816 2 3 4126 XOR2X2 $T=2025540 1874320 1 180 $X=2018940 $Y=1873918
X1088 8004 8002 2 3 3876 XOR2X2 $T=2067780 1894480 0 180 $X=2061180 $Y=1889040
X1089 8115 8111 2 3 4396 XOR2X2 $T=2098140 1834000 0 180 $X=2091540 $Y=1828560
X1090 9518 9505 2 3 779 XOR2X2 $T=2416920 1985200 0 180 $X=2410320 $Y=1979760
X1091 822 10095 2 3 818 XOR2X2 $T=2538360 1924720 0 180 $X=2531760 $Y=1919280
X1092 10271 10270 2 3 9492 XOR2X2 $T=2572020 1823920 1 180 $X=2565420 $Y=1823518
X1093 852 10433 2 3 9120 XOR2X2 $T=2611620 1813840 0 180 $X=2605020 $Y=1808400
X1094 2025 3 72 2 INVX2 $T=737220 1783600 1 0 $X=737218 $Y=1778160
X1095 155 3 218 2 INVX2 $T=1158960 1985200 0 0 $X=1158958 $Y=1984798
X1096 284 3 292 2 INVX2 $T=1305480 1924720 1 0 $X=1305478 $Y=1919280
X1097 5186 3 5210 2 INVX2 $T=1432200 1914640 0 180 $X=1430220 $Y=1909200
X1098 453 3 456 2 INVX2 $T=1614360 1874320 0 0 $X=1614358 $Y=1873918
X1099 611 3 7234 2 INVX2 $T=2055900 1924720 0 0 $X=2055898 $Y=1924318
X1100 557 3 6923 2 INVX2 $T=2108040 1924720 1 0 $X=2108038 $Y=1919280
X1101 8317 3 726 2 INVX2 $T=2220240 1985200 1 0 $X=2220238 $Y=1979760
X1102 8904 3 8930 2 INVX2 $T=2288220 1823920 1 0 $X=2288218 $Y=1818480
X1103 3522 2 3 3504 INVXL $T=1081080 1975120 1 180 $X=1079760 $Y=1974718
X1104 3463 2 3 3534 INVXL $T=1083060 1803760 0 0 $X=1083058 $Y=1803358
X1105 299 2 3 4746 INVXL $T=1340460 1834000 1 180 $X=1339140 $Y=1833598
X1106 4930 2 3 4901 INVXL $T=1374120 1954960 0 180 $X=1372800 $Y=1949520
X1107 5342 2 3 5324 INVXL $T=1461900 1904560 0 0 $X=1461898 $Y=1904158
X1108 5472 2 3 5467 INVXL $T=1487640 1914640 1 0 $X=1487638 $Y=1909200
X1109 5501 2 3 5560 INVXL $T=1500840 1914640 1 0 $X=1500838 $Y=1909200
X1110 139 2 3 419 INVXL $T=1544400 1834000 0 180 $X=1543080 $Y=1828560
X1111 5743 2 3 5721 INVXL $T=1552320 1914640 0 180 $X=1551000 $Y=1909200
X1112 5900 2 3 5917 INVXL $T=1592580 1894480 0 0 $X=1592578 $Y=1894078
X1113 541 2 3 6753 INVXL $T=1782660 1914640 1 180 $X=1781340 $Y=1914238
X1114 564 2 3 552 INVXL $T=1815000 1985200 0 0 $X=1814998 $Y=1984798
X1115 591 2 3 590 INVXL $T=1855920 1813840 0 180 $X=1854600 $Y=1808400
X1116 626 2 3 7838 INVXL $T=2026860 1834000 1 0 $X=2026858 $Y=1828560
X1117 603 2 3 8306 INVXL $T=2123880 1914640 0 0 $X=2123878 $Y=1914238
X1118 8444 2 3 8511 INVXL $T=2178660 1823920 0 0 $X=2178658 $Y=1823518
X1119 710 2 3 722 INVXL $T=2213640 1985200 1 180 $X=2212320 $Y=1984798
X1120 8978 2 3 9157 INVXL $T=2345640 1894480 1 180 $X=2344320 $Y=1894078
X1121 9072 2 3 9218 INVXL $T=2348280 1924720 0 0 $X=2348278 $Y=1924318
X1122 9044 2 3 9219 INVXL $T=2351580 1924720 0 0 $X=2351578 $Y=1924318
X1123 9023 2 3 9185 INVXL $T=2352900 1854160 0 180 $X=2351580 $Y=1848720
X1124 843 2 3 10405 INVXL $T=2597100 1783600 0 0 $X=2597098 $Y=1783198
X1125 4998 5102 4902 2 5030 5124 3 AOI31X1 $T=1405140 1934800 1 0 $X=1405138 $Y=1929360
X1126 5186 5523 5564 2 5565 5568 3 AOI31X1 $T=1502160 1924720 1 0 $X=1502158 $Y=1919280
X1127 10405 10409 853 2 858 10478 3 AOI31X1 $T=2620860 1793680 1 0 $X=2620858 $Y=1788240
X1128 2208 2271 2 3 2320 XNOR2X2 $T=785400 1924720 1 0 $X=785398 $Y=1919280
X1129 2381 2384 2 3 2498 XNOR2X2 $T=807840 1813840 0 0 $X=807838 $Y=1813438
X1130 2895 2900 2 3 3010 XNOR2X2 $T=931260 1823920 0 0 $X=931258 $Y=1823518
X1131 2948 2916 2 3 3058 XNOR2X2 $T=942480 1884400 1 0 $X=942478 $Y=1878960
X1132 7853 7921 2 3 4033 XNOR2X2 $T=2049300 1874320 0 180 $X=2042040 $Y=1868880
X1133 8057 8051 2 3 3918 XNOR2X2 $T=2081640 1864240 0 180 $X=2074380 $Y=1858800
X1134 676 675 2 3 7998 XNOR2X2 $T=2090880 1793680 0 180 $X=2083620 $Y=1788240
X1135 9453 9460 2 3 773 XNOR2X2 $T=2405700 1985200 0 180 $X=2398440 $Y=1979760
X1136 9573 9570 2 3 784 XNOR2X2 $T=2428800 1985200 0 180 $X=2421540 $Y=1979760
X1137 2362 2279 3 2 2369 XOR2X1 $T=799260 1934800 1 0 $X=799258 $Y=1929360
X1138 2405 98 3 2 2363 XOR2X1 $T=815100 1793680 0 180 $X=809820 $Y=1788240
X1139 99 100 3 2 2206 XOR2X1 $T=822360 1783600 0 180 $X=817080 $Y=1778160
X1140 101 2383 3 2 2448 XOR2X1 $T=820380 1954960 0 0 $X=820378 $Y=1954558
X1141 2511 2477 3 2 2491 XOR2X1 $T=844140 1844080 0 180 $X=838860 $Y=1838640
X1142 2709 2656 3 2 2841 XOR2X1 $T=885060 1874320 1 0 $X=885058 $Y=1868880
X1143 2805 2781 3 2 2806 XOR2X1 $T=904200 1854160 0 0 $X=904198 $Y=1853758
X1144 2820 2823 3 2 2842 XOR2X1 $T=909480 1904560 0 0 $X=909478 $Y=1904158
X1145 3098 3132 3 2 3152 XOR2X1 $T=985380 1854160 1 0 $X=985378 $Y=1848720
X1146 3211 3174 3 2 3241 XOR2X1 $T=1003200 1904560 0 0 $X=1003198 $Y=1904158
X1147 154 153 3 2 3212 XOR2X1 $T=1026960 1783600 0 180 $X=1021680 $Y=1778160
X1148 68 58 3 2 3293 XOR2X1 $T=1033560 1844080 0 180 $X=1028280 $Y=1838640
X1149 3338 156 3 2 3321 XOR2X1 $T=1040160 1783600 1 180 $X=1034880 $Y=1783198
X1150 3339 3417 3 2 3622 XOR2X1 $T=1052040 1874320 1 0 $X=1052038 $Y=1868880
X1151 3366 3437 3 2 3460 XOR2X1 $T=1058640 1904560 0 0 $X=1058638 $Y=1904158
X1152 180 179 3 2 3450 XOR2X1 $T=1071840 1975120 1 180 $X=1066560 $Y=1974718
X1153 3567 3566 3 2 3514 XOR2X1 $T=1089660 1823920 1 180 $X=1084380 $Y=1823518
X1154 3673 3711 3 2 3932 XOR2X1 $T=1118040 1914640 1 0 $X=1118038 $Y=1909200
X1155 3893 3892 3 2 3878 XOR2X1 $T=1157640 1904560 1 180 $X=1152360 $Y=1904158
X1156 3965 3962 3 2 217 XOR2X1 $T=1173480 1823920 0 180 $X=1168200 $Y=1818480
X1157 249 4240 3 2 3791 XOR2X1 $T=1228260 1934800 0 180 $X=1222980 $Y=1929360
X1158 4224 4264 3 2 4288 XOR2X1 $T=1229580 1894480 0 0 $X=1229578 $Y=1894078
X1159 260 4360 3 2 4202 XOR2X1 $T=1249380 1985200 0 180 $X=1244100 $Y=1979760
X1160 4408 4436 3 2 4453 XOR2X1 $T=1262580 1904560 1 0 $X=1262578 $Y=1899120
X1161 273 272 3 2 4449 XOR2X1 $T=1277100 1975120 1 180 $X=1271820 $Y=1974718
X1162 4456 276 3 2 3934 XOR2X1 $T=1278420 1934800 1 180 $X=1273140 $Y=1934398
X1163 4562 282 3 2 4503 XOR2X1 $T=1296900 1985200 0 180 $X=1291620 $Y=1979760
X1164 4611 4672 3 2 4694 XOR2X1 $T=1320000 1874320 0 0 $X=1319998 $Y=1873918
X1165 4687 4635 3 2 298 XOR2X1 $T=1323300 1803760 1 0 $X=1323298 $Y=1798320
X1166 304 4765 3 2 311 XOR2X1 $T=1341120 1823920 0 0 $X=1341118 $Y=1823518
X1167 4842 4750 3 2 315 XOR2X1 $T=1351680 1844080 0 0 $X=1351678 $Y=1843678
X1168 4914 4900 3 2 4918 XOR2X1 $T=1369500 1934800 0 0 $X=1369498 $Y=1934398
X1169 5010 5009 3 2 5028 XOR2X1 $T=1393260 1904560 0 0 $X=1393258 $Y=1904158
X1170 5084 5080 3 2 331 XOR2X1 $T=1404480 1854160 1 180 $X=1399200 $Y=1853758
X1171 5088 5083 3 2 337 XOR2X1 $T=1403820 1834000 0 0 $X=1403818 $Y=1833598
X1172 5126 5124 3 2 5088 XOR2X1 $T=1413060 1914640 1 180 $X=1407780 $Y=1914238
X1173 4863 5130 3 2 5121 XOR2X1 $T=1415700 1803760 0 180 $X=1410420 $Y=1798320
X1174 5227 5210 3 2 5084 XOR2X1 $T=1437480 1894480 0 180 $X=1432200 $Y=1889040
X1175 5269 5260 3 2 5235 XOR2X1 $T=1448040 1904560 1 180 $X=1442760 $Y=1904158
X1176 5713 5568 3 2 416 XOR2X1 $T=1539780 1874320 0 180 $X=1534500 $Y=1868880
X1177 5934 5931 3 2 440 XOR2X1 $T=1589940 1884400 0 180 $X=1584660 $Y=1878960
X1178 5951 5939 3 2 5934 XOR2X1 $T=1602480 1904560 0 180 $X=1597200 $Y=1899120
X1179 6349 6401 3 2 6377 XOR2X1 $T=1699500 1944880 1 180 $X=1694220 $Y=1944478
X1180 6782 6783 3 2 6681 XOR2X1 $T=1791900 1975120 0 180 $X=1786620 $Y=1969680
X1181 7586 7571 3 2 4395 XOR2X1 $T=1972740 1894480 0 180 $X=1967460 $Y=1889040
X1182 7566 7589 3 2 7468 XOR2X1 $T=1974060 1854160 1 180 $X=1968780 $Y=1853758
X1183 7644 7623 3 2 632 XOR2X1 $T=1984620 1975120 1 0 $X=1984618 $Y=1969680
X1184 7677 7676 3 2 7657 XOR2X1 $T=1995180 1854160 1 180 $X=1989900 $Y=1853758
X1185 473 618 3 2 7762 XOR2X1 $T=1994520 1823920 0 0 $X=1994518 $Y=1823518
X1186 639 7837 3 2 7781 XOR2X1 $T=2028840 1823920 0 180 $X=2023560 $Y=1818480
X1187 6983 607 3 2 7930 XOR2X1 $T=2040060 1924720 0 0 $X=2040058 $Y=1924318
X1188 7975 7981 3 2 7961 XOR2X1 $T=2060520 1823920 0 180 $X=2055240 $Y=1818480
X1189 8190 8183 3 2 686 XOR2X1 $T=2107380 1985200 0 0 $X=2107378 $Y=1984798
X1190 7098 607 3 2 8338 XOR2X1 $T=2120580 1894480 0 0 $X=2120578 $Y=1894078
X1191 7234 541 3 2 8411 XOR2X1 $T=2166120 1884400 0 180 $X=2160840 $Y=1878960
X1192 705 689 3 2 8445 XOR2X1 $T=2168760 1783600 0 0 $X=2168758 $Y=1783198
X1193 8585 8526 3 2 715 XOR2X1 $T=2204400 1823920 1 180 $X=2199120 $Y=1823518
X1194 8715 8716 3 2 8812 XOR2X1 $T=2238060 1965040 0 0 $X=2238058 $Y=1964638
X1195 8830 8835 3 2 8921 XOR2X1 $T=2267100 1975120 1 0 $X=2267098 $Y=1969680
X1196 9139 9114 3 2 9142 XOR2X1 $T=2337720 1944880 0 0 $X=2337718 $Y=1944478
X1197 781 780 3 2 9482 XOR2X1 $T=2413620 1803760 0 180 $X=2408340 $Y=1798320
X1198 788 8396 3 2 9650 XOR2X1 $T=2452560 1783600 1 180 $X=2447280 $Y=1783198
X1199 9780 9779 3 2 9269 XOR2X1 $T=2475000 1894480 1 180 $X=2469720 $Y=1894078
X1200 10263 10255 3 2 10214 XOR2X1 $T=2568060 1894480 0 180 $X=2562780 $Y=1889040
X1201 2451 2 2480 2528 3 NOR2BX1 $T=834240 1944880 1 0 $X=834238 $Y=1939440
X1202 114 2 53 117 3 NOR2BX1 $T=916080 1783600 1 0 $X=916078 $Y=1778160
X1203 3339 2 3416 3453 3 NOR2BX1 $T=1052040 1864240 1 0 $X=1052038 $Y=1858800
X1204 338 2 5167 5203 3 NOR2BX1 $T=1422960 1793680 0 0 $X=1422958 $Y=1793278
X1205 394 2 5499 5521 3 NOR2BX1 $T=1498200 1783600 1 0 $X=1498198 $Y=1778160
X1206 426 2 5860 5863 3 NOR2BX1 $T=1568160 1793680 0 0 $X=1568158 $Y=1793278
X1207 6222 2 6253 6256 3 NOR2BX1 $T=1661220 1965040 1 0 $X=1661218 $Y=1959600
X1208 7350 2 7317 4613 3 NOR2BX1 $T=1908720 1844080 1 180 $X=1906080 $Y=1843678
X1209 7384 2 7371 6442 3 NOR2BX1 $T=1927200 1954960 0 180 $X=1924560 $Y=1949520
X1210 8624 2 8596 8712 3 NOR2BX1 $T=2227500 1985200 1 0 $X=2227498 $Y=1979760
X1211 9922 2 806 9966 3 NOR2BX1 $T=2509980 1965040 1 0 $X=2509978 $Y=1959600
X1212 10099 2 729 10127 3 NOR2BX1 $T=2539020 1954960 1 0 $X=2539018 $Y=1949520
X1213 836 2 832 10325 3 NOR2BX1 $T=2583900 1944880 1 0 $X=2583898 $Y=1939440
X1214 46 31 36 28 2 3 1737 ADDFX2 $T=674520 1874320 0 180 $X=660660 $Y=1868880
X1215 21 1737 1769 44 2 3 1874 ADDFX2 $T=661320 1854160 0 0 $X=661318 $Y=1853758
X1216 50 46 22 37 2 3 34 ADDFX2 $T=678480 1834000 1 180 $X=664620 $Y=1833598
X1217 53 49 45 43 2 3 40 ADDFX2 $T=682440 1803760 0 180 $X=668580 $Y=1798320
X1218 62 53 49 52 2 3 48 ADDFX2 $T=690360 1894480 1 180 $X=676500 $Y=1894078
X1219 1795 1807 1826 1835 2 3 1850 ADDFX2 $T=679800 1854160 1 0 $X=679798 $Y=1848720
X1220 58 55 36 24 2 3 51 ADDFX2 $T=693660 1934800 1 180 $X=679800 $Y=1934398
X1221 49 55 58 1842 2 3 1795 ADDFX2 $T=681120 1884400 1 0 $X=681118 $Y=1878960
X1222 36 42 45 1810 2 3 1807 ADDFX2 $T=696300 1844080 0 180 $X=682440 $Y=1838640
X1223 1842 1841 1810 54 2 3 1796 ADDFX2 $T=696960 1874320 1 180 $X=683100 $Y=1873918
X1224 41 36 45 1870 2 3 1947 ADDFX2 $T=687720 1944880 1 0 $X=687718 $Y=1939440
X1225 57 31 1870 1826 2 3 1930 ADDFX2 $T=689040 1914640 1 0 $X=689038 $Y=1909200
X1226 53 58 55 1931 2 3 63 ADDFX2 $T=722040 1985200 1 180 $X=708180 $Y=1984798
X1227 55 46 1841 1986 2 3 1969 ADDFX2 $T=710160 1884400 0 0 $X=710158 $Y=1883998
X1228 49 23 22 2054 2 3 2074 ADDFX2 $T=737880 1894480 1 0 $X=737878 $Y=1889040
X1229 2091 2074 1986 2029 2 3 1968 ADDFX2 $T=751740 1884400 0 180 $X=737880 $Y=1878960
X1230 62 53 46 2030 2 3 2091 ADDFX2 $T=762300 1864240 1 180 $X=748440 $Y=1863838
X1231 53 46 104 2476 2 3 2499 ADDFX2 $T=826320 1985200 0 0 $X=826318 $Y=1984798
X1232 108 109 110 2591 2 3 2589 ADDFX2 $T=850080 1793680 0 0 $X=850078 $Y=1793278
X1233 62 55 50 2614 2 3 2732 ADDFX2 $T=902880 1944880 1 180 $X=889020 $Y=1944478
X1234 345 319 349 5234 2 3 5214 ADDFX2 $T=1427580 1985200 0 0 $X=1427578 $Y=1984798
X1235 430 238 422 5765 2 3 5746 ADDFX2 $T=1560240 1985200 0 180 $X=1546380 $Y=1979760
X1236 308 428 354 5839 2 3 5821 ADDFX2 $T=1552980 1944880 0 0 $X=1552978 $Y=1944478
X1237 435 418 429 5805 2 3 5772 ADDFX2 $T=1566840 1975120 1 180 $X=1552980 $Y=1974718
X1238 6218 469 6161 6152 2 3 466 ADDFX2 $T=1654620 1934800 0 180 $X=1640760 $Y=1929360
X1239 7420 7425 7416 7401 2 3 4733 ADDFX2 $T=1945680 1874320 0 180 $X=1931820 $Y=1868880
X1240 7407 582 607 7776 2 3 7699 ADDFX2 $T=2021580 1944880 0 180 $X=2007720 $Y=1939440
X1241 7234 6923 7857 7840 2 3 7783 ADDFX2 $T=2041380 1965040 0 180 $X=2027520 $Y=1959600
X1242 7930 6811 7897 7881 2 3 7879 ADDFX2 $T=2050620 1944880 0 180 $X=2036760 $Y=1939440
X1243 8094 7234 8059 8052 2 3 8039 ADDFX2 $T=2090220 1954960 0 180 $X=2076360 $Y=1949520
X1244 8167 6923 8087 8096 2 3 8091 ADDFX2 $T=2104080 1944880 1 180 $X=2090220 $Y=1944478
X1245 7032 603 702 8469 2 3 8540 ADDFX2 $T=2166120 1934800 0 0 $X=2166118 $Y=1934398
X1246 6983 559 6751 8474 2 3 8537 ADDFX2 $T=2170740 1914640 0 0 $X=2170738 $Y=1914238
X1247 6751 606 6923 8475 2 3 8616 ADDFX2 $T=2170740 1954960 0 0 $X=2170738 $Y=1954558
X1248 713 575 541 8598 2 3 8601 ADDFX2 $T=2194500 1914640 1 0 $X=2194498 $Y=1909200
X1249 7098 582 719 8621 2 3 8641 ADDFX2 $T=2200440 1904560 1 0 $X=2200438 $Y=1899120
X1250 611 725 6811 8676 2 3 8743 ADDFX2 $T=2216280 1934800 1 0 $X=2216278 $Y=1929360
X1251 8705 718 8774 8779 2 3 8939 ADDFX2 $T=2242020 1834000 0 0 $X=2242018 $Y=1833598
X1252 709 530 8816 736 2 3 8831 ADDFX2 $T=2254560 1793680 0 0 $X=2254558 $Y=1793278
X1253 2090 2092 3 2 79 XNOR2X1 $T=747780 1924720 1 0 $X=747778 $Y=1919280
X1254 1975 1998 3 2 2134 XNOR2X1 $T=749760 1823920 1 0 $X=749758 $Y=1818480
X1255 2194 2154 3 2 2211 XNOR2X1 $T=768240 1934800 1 0 $X=768238 $Y=1929360
X1256 2479 2478 3 2 2367 XNOR2X1 $T=836220 1834000 1 180 $X=830940 $Y=1833598
X1257 2528 2529 3 2 2613 XNOR2X1 $T=847440 1924720 0 0 $X=847438 $Y=1924318
X1258 2527 2653 3 2 2840 XNOR2X1 $T=870540 1864240 1 0 $X=870538 $Y=1858800
X1259 2703 2724 3 2 2700 XNOR2X1 $T=885720 1844080 0 0 $X=885718 $Y=1843678
X1260 2780 2697 3 2 2938 XNOR2X1 $T=912780 1894480 1 0 $X=912778 $Y=1889040
X1261 112 3142 3 2 3106 XNOR2X1 $T=990660 1834000 0 180 $X=985380 $Y=1828560
X1262 150 3224 3 2 3114 XNOR2X1 $T=1006500 1844080 0 180 $X=1001220 $Y=1838640
X1263 3138 3225 3 2 3513 XNOR2X1 $T=1003860 1894480 0 0 $X=1003858 $Y=1894078
X1264 3137 3258 3 2 3475 XNOR2X1 $T=1016400 1884400 1 0 $X=1016398 $Y=1878960
X1265 152 109 3 2 3299 XNOR2X1 $T=1026960 1813840 0 0 $X=1026958 $Y=1813438
X1266 3322 3358 3 2 3431 XNOR2X1 $T=1045440 1914640 0 0 $X=1045438 $Y=1914238
X1267 3480 3479 3 2 3457 XNOR2X1 $T=1068540 1783600 1 180 $X=1063260 $Y=1783198
X1268 3495 3547 3 2 3589 XNOR2X1 $T=1085040 1914640 1 0 $X=1085038 $Y=1909200
X1269 3610 3615 3 2 3592 XNOR2X1 $T=1100220 1834000 1 180 $X=1094940 $Y=1833598
X1270 3735 3656 3 2 3832 XNOR2X1 $T=1123980 1894480 0 0 $X=1123978 $Y=1894078
X1271 3811 3810 3 2 213 XNOR2X1 $T=1145100 1823920 1 180 $X=1139820 $Y=1823518
X1272 3749 3814 3 2 3933 XNOR2X1 $T=1145100 1864240 1 0 $X=1145098 $Y=1858800
X1273 3917 3914 3 2 3931 XNOR2X1 $T=1160940 1904560 1 0 $X=1160938 $Y=1899120
X1274 4125 4143 3 2 4178 XNOR2X1 $T=1207800 1904560 1 0 $X=1207798 $Y=1899120
X1275 4199 246 3 2 4030 XNOR2X1 $T=1218360 1944880 0 180 $X=1213080 $Y=1939440
X1276 4313 4348 3 2 4393 XNOR2X1 $T=1246740 1904560 1 0 $X=1246738 $Y=1899120
X1277 269 4457 3 2 4327 XNOR2X1 $T=1270500 1985200 1 180 $X=1265220 $Y=1984798
X1278 4471 4470 3 2 4431 XNOR2X1 $T=1273140 1823920 0 180 $X=1267860 $Y=1818480
X1279 279 4511 3 2 4495 XNOR2X1 $T=1283700 1924720 0 180 $X=1278420 $Y=1919280
X1280 4486 4539 3 2 4532 XNOR2X1 $T=1288980 1894480 1 0 $X=1288978 $Y=1889040
X1281 294 296 3 2 4684 XNOR2X1 $T=1316040 1975120 0 0 $X=1316038 $Y=1974718
X1282 299 4706 3 2 4668 XNOR2X1 $T=1330560 1834000 1 180 $X=1325280 $Y=1833598
X1283 313 314 3 2 4842 XNOR2X1 $T=1351680 1975120 1 0 $X=1351678 $Y=1969680
X1284 4918 4920 3 2 320 XNOR2X1 $T=1374780 1823920 0 180 $X=1369500 $Y=1818480
X1285 4928 4917 3 2 324 XNOR2X1 $T=1374120 1834000 1 0 $X=1374118 $Y=1828560
X1286 4949 4902 3 2 4921 XNOR2X1 $T=1375440 1934800 1 0 $X=1375438 $Y=1929360
X1287 5028 5027 3 2 330 XNOR2X1 $T=1398540 1844080 1 180 $X=1393260 $Y=1843678
X1288 5188 5204 3 2 351 XNOR2X1 $T=1432200 1894480 0 0 $X=1432198 $Y=1894078
X1289 5360 5359 3 2 361 XNOR2X1 $T=1463880 1904560 0 180 $X=1458600 $Y=1899120
X1290 5425 5424 3 2 376 XNOR2X1 $T=1479720 1904560 0 180 $X=1474440 $Y=1899120
X1291 5477 5471 3 2 388 XNOR2X1 $T=1488960 1874320 0 0 $X=1488958 $Y=1873918
X1292 5563 5567 3 2 396 XNOR2X1 $T=1506120 1884400 0 180 $X=1500840 $Y=1878960
X1293 5631 5632 3 2 404 XNOR2X1 $T=1520640 1874320 0 180 $X=1515360 $Y=1868880
X1294 5700 5696 3 2 413 XNOR2X1 $T=1538460 1894480 0 180 $X=1533180 $Y=1889040
X1295 418 417 3 2 415 XNOR2X1 $T=1539780 1985200 0 180 $X=1534500 $Y=1979760
X1296 5877 5875 3 2 436 XNOR2X1 $T=1574100 1864240 1 180 $X=1568820 $Y=1863838
X1297 6135 6133 3 2 6161 XNOR2X1 $T=1639440 1965040 1 0 $X=1639438 $Y=1959600
X1298 6304 6315 3 2 6326 XNOR2X1 $T=1675740 1954960 1 0 $X=1675738 $Y=1949520
X1299 6482 6502 3 2 6518 XNOR2X1 $T=1717980 1954960 1 0 $X=1717978 $Y=1949520
X1300 7173 603 3 2 6083 XNOR2X1 $T=1877040 1975120 1 180 $X=1871760 $Y=1974718
X1301 7401 7417 3 2 4550 XNOR2X1 $T=1938420 1894480 0 180 $X=1933140 $Y=1889040
X1302 7407 603 3 2 7420 XNOR2X1 $T=1934460 1924720 0 0 $X=1934458 $Y=1924318
X1303 7440 7426 3 2 7372 XNOR2X1 $T=1942380 1954960 1 180 $X=1937100 $Y=1954558
X1304 7445 7526 3 2 4489 XNOR2X1 $T=1960860 1894480 1 180 $X=1955580 $Y=1894078
X1305 626 625 3 2 7439 XNOR2X1 $T=1963500 1844080 1 180 $X=1958220 $Y=1843678
X1306 7636 7637 3 2 4312 XNOR2X1 $T=1984620 1874320 0 180 $X=1979340 $Y=1868880
X1307 7761 7821 3 2 7683 XNOR2X1 $T=2026200 1844080 1 180 $X=2020920 $Y=1843678
X1308 7924 7923 3 2 7864 XNOR2X1 $T=2049960 1793680 1 180 $X=2044680 $Y=1793278
X1309 639 625 3 2 8213 XNOR2X1 $T=2107380 1783600 1 0 $X=2107378 $Y=1778160
X1310 8393 8391 3 2 699 XNOR2X1 $T=2155560 1834000 0 180 $X=2150280 $Y=1828560
X1311 8496 708 3 2 8443 XNOR2X1 $T=2188560 1834000 0 180 $X=2183280 $Y=1828560
X1312 725 557 3 2 8672 XNOR2X1 $T=2220900 1904560 0 0 $X=2220898 $Y=1904158
X1313 725 6753 3 2 8710 XNOR2X1 $T=2230140 1854160 0 0 $X=2230138 $Y=1853758
X1314 729 550 3 2 8774 XNOR2X1 $T=2243340 1813840 1 0 $X=2243338 $Y=1808400
X1315 732 8622 3 2 731 XNOR2X1 $T=2248620 1823920 0 180 $X=2243340 $Y=1818480
X1316 713 532 3 2 8772 XNOR2X1 $T=2244660 1874320 0 0 $X=2244658 $Y=1873918
X1317 9105 9108 3 2 9241 XNOR2X1 $T=2329800 1954960 0 0 $X=2329798 $Y=1954558
X1318 9111 9093 3 2 9137 XNOR2X1 $T=2332440 1844080 1 0 $X=2332438 $Y=1838640
X1319 9033 9173 3 2 9167 XNOR2X1 $T=2343000 1823920 0 0 $X=2342998 $Y=1823518
X1320 9227 9222 3 2 9274 XNOR2X1 $T=2355540 1904560 1 0 $X=2355538 $Y=1899120
X1321 9220 9235 3 2 9316 XNOR2X1 $T=2355540 1954960 1 0 $X=2355538 $Y=1949520
X1322 9272 9273 3 2 9458 XNOR2X1 $T=2368080 1874320 1 0 $X=2368078 $Y=1868880
X1323 8942 9286 3 2 9477 XNOR2X1 $T=2370060 1904560 1 0 $X=2370058 $Y=1899120
X1324 9304 9307 3 2 9459 XNOR2X1 $T=2375340 1914640 1 0 $X=2375338 $Y=1909200
X1325 9482 9484 3 2 9497 XNOR2X1 $T=2407020 1813840 1 0 $X=2407018 $Y=1808400
X1326 9650 787 3 2 9706 XNOR2X1 $T=2447280 1793680 0 0 $X=2447278 $Y=1793278
X1327 729 10099 3 2 10148 XNOR2X1 $T=2537700 1965040 1 0 $X=2537698 $Y=1959600
X1328 3877 3809 3 108 2 215 3794 214 OAI221XL $T=1145100 1783600 1 180 $X=1140480 $Y=1783198
X1329 5342 5258 3 5210 2 5343 5321 5360 OAI221XL $T=1459260 1914640 0 0 $X=1459258 $Y=1914238
X1330 5472 5426 3 5210 2 5478 5442 5471 OAI221XL $T=1492260 1904560 1 180 $X=1487640 $Y=1904158
X1331 5588 5210 3 5426 2 5560 5559 5567 OAI221XL $T=1508100 1904560 1 180 $X=1503480 $Y=1904158
X1332 5800 5846 3 5838 2 5841 5862 5900 OAI221XL $T=1566180 1894480 0 0 $X=1566178 $Y=1894078
X1333 7097 7099 3 575 2 7014 7008 7048 OAI221XL $T=1850640 1844080 1 180 $X=1846020 $Y=1843678
X1334 8993 8995 3 9029 2 8977 9028 9025 OAI221XL $T=2311980 1854160 1 0 $X=2311978 $Y=1848720
X1335 8993 9185 3 9090 2 9163 8977 9168 OAI221XL $T=2344980 1854160 0 180 $X=2340360 $Y=1848720
X1336 10253 10065 3 10254 2 10252 10053 10215 OAI221XL $T=2567400 1934800 0 180 $X=2562780 $Y=1929360
X1337 112 2636 111 2 3 2586 ADDHXL $T=870540 1834000 0 180 $X=863280 $Y=1828560
X1338 5208 5165 333 2 3 5130 ADDHXL $T=1435500 1803760 0 180 $X=1428240 $Y=1798320
X1339 5320 5274 358 2 3 5208 ADDHXL $T=1455960 1803760 0 180 $X=1448700 $Y=1798320
X1340 5364 364 363 2 3 5320 ADDHXL $T=1466520 1793680 0 180 $X=1459260 $Y=1788240
X1341 383 5447 381 2 3 5364 ADDHXL $T=1488960 1783600 0 180 $X=1481700 $Y=1778160
X1342 303 5921 428 2 3 5975 ADDHXL $T=1582020 1934800 0 0 $X=1582018 $Y=1934398
X1343 6015 6014 148 2 3 438 ADDHXL $T=1605780 1783600 0 180 $X=1598520 $Y=1778160
X1344 467 6142 149 2 3 6015 ADDHXL $T=1646700 1783600 0 180 $X=1639440 $Y=1778160
X1345 6983 7591 7305 2 3 7679 ADDHXL $T=1987260 1934800 0 0 $X=1987258 $Y=1934398
X1346 7032 7857 7305 2 3 7897 ADDHXL $T=2029500 1934800 0 0 $X=2029498 $Y=1934398
X1347 541 8059 7032 2 3 8087 ADDHXL $T=2077020 1944880 0 0 $X=2077018 $Y=1944478
X1348 6751 8326 8306 2 3 8313 ADDHXL $T=2146320 1914640 1 180 $X=2139060 $Y=1914238
X1349 2 62 111 3416 3 NOR2XL $T=1052040 1854160 1 0 $X=1052038 $Y=1848720
X1350 2 180 173 3477 3 NOR2XL $T=1063920 1965040 0 0 $X=1063918 $Y=1964638
X1351 2 185 192 3515 3 NOR2XL $T=1089660 1803760 0 180 $X=1087680 $Y=1798320
X1352 2 272 273 4457 3 NOR2XL $T=1277760 1985200 1 180 $X=1275780 $Y=1984798
X1353 2 276 4456 4511 3 NOR2XL $T=1279740 1934800 1 0 $X=1279738 $Y=1929360
X1354 2 5692 5715 5799 3 NOR2XL $T=1555620 1914640 1 0 $X=1555618 $Y=1909200
X1355 2 319 5975 5988 3 NOR2XL $T=1613040 1934800 1 180 $X=1611060 $Y=1934398
X1356 2 6239 472 6253 3 NOR2XL $T=1660560 1975120 1 0 $X=1660558 $Y=1969680
X1357 2 559 7367 7317 3 NOR2XL $T=1922580 1844080 1 180 $X=1920600 $Y=1843678
X1358 2 7367 7372 7371 3 NOR2XL $T=1926540 1944880 0 180 $X=1924560 $Y=1939440
X1359 2 626 639 7996 3 NOR2XL $T=2060520 1834000 0 0 $X=2060518 $Y=1833598
X1360 2 575 606 8094 3 NOR2XL $T=2086920 1965040 0 0 $X=2086918 $Y=1964638
X1361 2 8983 9138 9129 3 NOR2XL $T=2339700 1864240 1 180 $X=2337720 $Y=1863838
X1362 81 84 87 3 2 2291 XOR3X2 $T=804540 1985200 1 180 $X=792660 $Y=1984798
X1363 2695 2750 2732 3 2 2772 XOR3X2 $T=909480 1934800 0 180 $X=897600 $Y=1929360
X1364 155 160 3357 3 2 167 XOR3X2 $T=1034880 1823920 0 0 $X=1034878 $Y=1823518
X1365 3429 168 164 3 2 162 XOR3X2 $T=1055340 1803760 0 180 $X=1043460 $Y=1798320
X1366 3543 188 186 3 2 184 XOR3X2 $T=1083720 1954960 0 180 $X=1071840 $Y=1949520
X1367 193 190 3521 3 2 189 XOR3X2 $T=1089000 1864240 1 180 $X=1077120 $Y=1863838
X1368 211 205 3689 3 2 203 XOR3X2 $T=1122000 1834000 1 180 $X=1110120 $Y=1833598
X1369 5766 5765 5772 3 2 431 XOR3X2 $T=1549020 1914640 0 0 $X=1549018 $Y=1914238
X1370 5771 5805 5821 3 2 432 XOR3X2 $T=1549680 1874320 1 0 $X=1549678 $Y=1868880
X1371 5901 5932 5921 3 2 444 XOR3X2 $T=1581360 1914640 0 0 $X=1581358 $Y=1914238
X1372 5964 417 319 3 2 439 XOR3X2 $T=1595880 1944880 0 180 $X=1584000 $Y=1939440
X1373 7610 7591 7234 3 2 7543 XOR3X2 $T=1981320 1934800 1 180 $X=1969440 $Y=1934398
X1374 638 7783 7776 3 2 641 XOR3X2 $T=2008380 1985200 0 0 $X=2008378 $Y=1984798
X1375 759 9162 757 3 2 755 XOR3X2 $T=2349600 1783600 0 180 $X=2337720 $Y=1778160
X1376 9325 9280 764 3 2 763 XOR3X2 $T=2377320 1823920 0 180 $X=2365440 $Y=1818480
X1377 9538 9498 9486 3 2 9042 XOR3X2 $T=2419560 1864240 0 180 $X=2407680 $Y=1858800
X1378 9615 9708 9707 3 2 9156 XOR3X2 $T=2460480 1874320 1 180 $X=2448600 $Y=1873918
X1379 789 9744 793 3 2 9707 XOR3X2 $T=2458500 1803760 0 0 $X=2458498 $Y=1803358
X1380 797 798 800 3 2 9811 XOR3X2 $T=2484900 1803760 1 0 $X=2484898 $Y=1798320
X1381 9865 9836 9831 3 2 9318 XOR3X2 $T=2496780 1884400 0 180 $X=2484900 $Y=1878960
X1382 10216 828 10082 3 2 9576 XOR3X2 $T=2554200 1834000 0 180 $X=2542320 $Y=1828560
X1383 5561 5428 2 5566 3 5569 AOI21XL $T=1502820 1944880 1 0 $X=1502818 $Y=1939440
X1384 5605 5615 2 5606 3 5629 AOI21XL $T=1515360 1904560 0 0 $X=1515358 $Y=1904158
X1385 9000 9073 2 9021 3 9135 AOI21XL $T=2325840 1884400 1 0 $X=2325838 $Y=1878960
X1386 9219 9040 2 9218 3 9270 AOI21XL $T=2356860 1924720 0 0 $X=2356858 $Y=1924318
X1387 2154 2067 2136 3 2092 2 OAI2BB1X1 $T=753720 1934800 0 180 $X=750420 $Y=1929360
X1388 2401 95 2299 3 2384 2 OAI2BB1X1 $T=811800 1834000 0 180 $X=808500 $Y=1828560
X1389 196 3564 193 3 3542 2 OAI2BB1X1 $T=1091640 1884400 0 180 $X=1088340 $Y=1878960
X1390 3749 3738 3734 3 3735 2 OAI2BB1X1 $T=1127940 1864240 1 180 $X=1124640 $Y=1863838
X1391 219 235 4073 3 4121 2 OAI2BB1X1 $T=1199220 1783600 1 0 $X=1199218 $Y=1778160
X1392 5252 5186 5258 3 5260 2 OAI2BB1X1 $T=1444080 1914640 0 0 $X=1444078 $Y=1914238
X1393 6135 6080 6129 3 6304 2 OAI2BB1X1 $T=1638780 1975120 1 0 $X=1638778 $Y=1969680
X1394 572 6877 584 3 7002 2 OAI2BB1X1 $T=1837440 1803760 1 0 $X=1837438 $Y=1798320
X1395 7401 7406 7403 3 7445 2 OAI2BB1X1 $T=1937100 1894480 0 0 $X=1937098 $Y=1894078
X1396 7470 7426 7472 3 7610 2 OAI2BB1X1 $T=1954260 1954960 0 0 $X=1954258 $Y=1954558
X1397 7995 7960 7974 3 7923 2 OAI2BB1X1 $T=2061840 1793680 1 180 $X=2058540 $Y=1793278
X1398 8679 8602 8595 3 8717 2 OAI2BB1X1 $T=2230140 1975120 1 0 $X=2230138 $Y=1969680
X1399 8624 726 8782 3 8796 2 OAI2BB1X1 $T=2251920 1985200 1 0 $X=2251918 $Y=1979760
X1400 9073 9027 9039 3 9019 2 OAI2BB1X1 $T=2317260 1874320 0 180 $X=2313960 $Y=1868880
X1401 9084 8659 9076 3 9093 2 OAI2BB1X1 $T=2326500 1874320 0 0 $X=2326498 $Y=1873918
X1402 9026 8659 9116 3 9222 2 OAI2BB1X1 $T=2350260 1904560 1 0 $X=2350258 $Y=1899120
X1403 775 782 783 3 9543 2 OAI2BB1X1 $T=2415600 1783600 1 0 $X=2415598 $Y=1778160
X1404 9376 9504 9494 3 9498 2 OAI2BB1X1 $T=2420220 1854160 1 180 $X=2416920 $Y=1853758
X1405 781 9484 9525 3 9486 2 OAI2BB1X1 $T=2418900 1803760 0 0 $X=2418898 $Y=1803358
X1406 788 787 8396 3 9724 2 OAI2BB1X1 $T=2455860 1783600 0 0 $X=2455858 $Y=1783198
X1407 9722 786 9723 3 9708 2 OAI2BB1X1 $T=2458500 1854160 1 0 $X=2458498 $Y=1848720
X1408 789 793 9745 3 9759 2 OAI2BB1X1 $T=2463780 1823920 1 0 $X=2463778 $Y=1818480
X1409 797 800 9837 3 9831 2 OAI2BB1X1 $T=2493480 1793680 0 180 $X=2490180 $Y=1788240
X1410 817 823 10152 3 10216 2 OAI2BB1X1 $T=2547600 1803760 0 0 $X=2547598 $Y=1803358
X1411 10321 837 841 3 10320 2 OAI2BB1X1 $T=2583900 1954960 1 0 $X=2583898 $Y=1949520
X1412 10405 10412 845 3 10465 2 OAI2BB1X1 $T=2614260 1783600 0 0 $X=2614258 $Y=1783198
X1413 10465 853 10478 3 859 2 OAI2BB1X1 $T=2620200 1783600 0 0 $X=2620198 $Y=1783198
X1414 1997 3 2050 2 74 NAND2BXL $T=749760 1803760 1 180 $X=747120 $Y=1803358
X1415 114 3 53 2 116 NAND2BXL $T=900240 1783600 1 180 $X=897600 $Y=1783198
X1416 210 3 112 2 3795 NAND2BXL $T=1139820 1803760 0 0 $X=1139818 $Y=1803358
X1417 3873 3 3820 2 3801 NAND2BXL $T=1147740 1874320 0 180 $X=1145100 $Y=1868880
X1418 4128 3 4079 2 4144 NAND2BXL $T=1205160 1864240 1 0 $X=1205158 $Y=1858800
X1419 4311 3 4286 2 3965 NAND2BXL $T=1236180 1823920 0 180 $X=1233540 $Y=1818480
X1420 4364 3 4339 2 4332 NAND2BXL $T=1246740 1864240 0 180 $X=1244100 $Y=1858800
X1421 4527 3 4516 2 4519 NAND2BXL $T=1290300 1864240 0 0 $X=1290298 $Y=1863838
X1422 4650 3 4649 2 4633 NAND2BXL $T=1314720 1844080 1 180 $X=1312080 $Y=1843678
X1423 5089 3 5122 2 5126 NAND2BXL $T=1417020 1965040 1 0 $X=1417018 $Y=1959600
X1424 5212 3 5213 2 5227 NAND2BXL $T=1435500 1904560 0 0 $X=1435498 $Y=1904158
X1425 5609 3 5610 2 5631 NAND2BXL $T=1523940 1954960 0 180 $X=1521300 $Y=1949520
X1426 521 3 500 2 6800 NAND2BXL $T=1791900 1823920 0 0 $X=1791898 $Y=1823518
X1427 582 3 574 2 7008 NAND2BXL $T=1838100 1854160 1 0 $X=1838098 $Y=1848720
X1428 8314 3 8316 2 697 NAND2BXL $T=2141700 1965040 0 0 $X=2141698 $Y=1964638
X1429 8504 3 8505 2 720 NAND2BXL $T=2188560 1985200 0 0 $X=2188558 $Y=1984798
X1430 8600 3 8639 2 8715 NAND2BXL $T=2223540 1965040 1 0 $X=2223538 $Y=1959600
X1431 8596 3 8595 2 8830 NAND2BXL $T=2253900 1975120 1 0 $X=2253898 $Y=1969680
X1432 8905 3 8919 2 8942 NAND2BXL $T=2290200 1884400 0 0 $X=2290198 $Y=1883998
X1433 9032 3 9041 2 9105 NAND2BXL $T=2319240 1954960 1 0 $X=2319238 $Y=1949520
X1434 8992 3 8887 2 9139 NAND2BXL $T=2332440 1944880 1 0 $X=2332438 $Y=1939440
X1435 10065 3 10053 2 10054 NAND2BXL $T=2528460 1934800 0 180 $X=2525820 $Y=1929360
X1436 1930 1948 1968 1975 2 3 1989 ADDFHX1 $T=706860 1874320 0 0 $X=706858 $Y=1873918
X1437 1931 1947 1969 1948 2 3 1965 ADDFHX1 $T=706860 1934800 0 0 $X=706858 $Y=1934398
X1438 64 67 1965 1972 2 3 2052 ADDFHX1 $T=706860 1975120 1 0 $X=706858 $Y=1969680
X1439 41 2030 2054 1769 2 3 2072 ADDFHX1 $T=726660 1854160 0 0 $X=726658 $Y=1853758
X1440 81 84 87 2195 2 3 2216 ADDFHX1 $T=759660 1985200 0 0 $X=759658 $Y=1984798
X1441 91 93 96 2275 2 3 2383 ADDFHX1 $T=785400 1985200 1 0 $X=785398 $Y=1979760
X1442 1757 3 39 2 1761 38 NAND3X1 $T=668580 1914640 1 180 $X=665940 $Y=1914238
X1443 418 417 319 5932 3 2 5951 CMPR32X1 $T=1580700 1965040 1 0 $X=1580698 $Y=1959600
X1444 310 377 450 5939 3 2 5864 CMPR32X1 $T=1618320 1965040 0 180 $X=1604460 $Y=1959600
X1445 2499 2614 2475 2634 2639 3 2 OAI2BB2X2 $T=862620 1954960 1 0 $X=862618 $Y=1949520
X1446 9972 9999 10064 3 10000 2 AOI2BB1X2 $T=2517240 1874320 1 0 $X=2517238 $Y=1868880
X1447 1796 1835 1874 1845 2 3 1912 ADDFHX2 $T=679140 1823920 0 0 $X=679138 $Y=1823518
X1448 2072 2029 1850 1963 2 3 1998 ADDFHX2 $T=747780 1834000 1 180 $X=725340 $Y=1833598
X1449 650 7878 3 2 7817 OR2X1 $T=2047320 1803760 0 180 $X=2044680 $Y=1798320
X1450 659 661 3 2 7976 OR2X1 $T=2055900 1864240 1 0 $X=2055898 $Y=1858800
X1451 95 2 2280 3 CLKINVX3 $T=788700 1834000 0 180 $X=786720 $Y=1828560
X1452 2475 2 2529 3 CLKINVX3 $T=846780 1954960 1 0 $X=846778 $Y=1949520
X1453 2878 2 2911 3 CLKINVX3 $T=927960 1813840 1 0 $X=927958 $Y=1808400
X1454 3292 2 3137 3 CLKINVX3 $T=1026300 1904560 0 180 $X=1024320 $Y=1899120
X1455 3546 2 3465 3 CLKINVX3 $T=1068540 1854160 0 180 $X=1066560 $Y=1848720
X1456 185 2 177 3 CLKINVX3 $T=1072500 1823920 0 0 $X=1072498 $Y=1823518
X1457 3715 2 3712 3 CLKINVX3 $T=1118700 1934800 0 0 $X=1118698 $Y=1934398
X1458 225 2 171 3 CLKINVX3 $T=1197240 1975120 1 0 $X=1197238 $Y=1969680
X1459 4843 2 317 3 CLKINVX3 $T=1357620 1874320 0 0 $X=1357618 $Y=1873918
X1460 377 2 319 3 CLKINVX3 $T=1471140 1975120 0 180 $X=1469160 $Y=1969680
X1461 5439 2 378 3 CLKINVX3 $T=1473780 1783600 0 180 $X=1471800 $Y=1778160
X1462 449 2 5973 3 CLKINVX3 $T=1603140 1864240 1 0 $X=1603138 $Y=1858800
X1463 451 2 452 3 CLKINVX3 $T=1611060 1894480 1 0 $X=1611058 $Y=1889040
X1464 459 2 460 3 CLKINVX3 $T=1628880 1904560 1 0 $X=1628878 $Y=1899120
X1465 511 2 6659 3 CLKINVX3 $T=1752960 1965040 1 0 $X=1752958 $Y=1959600
X1466 6779 2 541 3 CLKINVX3 $T=1787940 1904560 0 180 $X=1785960 $Y=1899120
X1467 6983 2 575 3 CLKINVX3 $T=1832820 1864240 0 0 $X=1832818 $Y=1863838
X1468 7119 2 7032 3 CLKINVX3 $T=1855920 1924720 0 0 $X=1855918 $Y=1924318
X1469 606 2 607 3 CLKINVX3 $T=1919280 1944880 1 0 $X=1919278 $Y=1939440
X1470 532 2 6811 3 CLKINVX3 $T=2068440 1914640 1 0 $X=2068438 $Y=1909200
X1471 707 2 702 3 CLKINVX3 $T=2180640 1854160 0 0 $X=2180638 $Y=1853758
X1472 619 2 589 3 CLKINVX3 $T=2209680 1844080 1 0 $X=2209678 $Y=1838640
X1473 724 2 709 3 CLKINVX3 $T=2224860 1783600 0 0 $X=2224858 $Y=1783198
X1474 713 2 738 3 CLKINVX3 $T=2269740 1823920 0 180 $X=2267760 $Y=1818480
X1475 9116 2 9073 3 CLKINVX3 $T=2337720 1904560 1 0 $X=2337718 $Y=1899120
X1476 8659 2 9114 3 CLKINVX3 $T=2347620 1934800 0 180 $X=2345640 $Y=1929360
X1477 164 168 2 3 3413 AND2X1 $T=1048080 1803760 0 0 $X=1048078 $Y=1803358
X1478 4474 3897 2 3 4485 AND2X1 $T=1273140 1854160 0 0 $X=1273138 $Y=1853758
X1479 4609 4611 2 3 4612 AND2X1 $T=1301520 1864240 0 0 $X=1301518 $Y=1863838
X1480 5324 5321 2 3 5269 AND2X1 $T=1454640 1904560 1 180 $X=1452000 $Y=1904158
X1481 6249 474 2 3 6251 AND2X1 $T=1661220 1834000 1 0 $X=1661218 $Y=1828560
X1482 7591 7234 2 3 7619 AND2X1 $T=1985940 1954960 1 0 $X=1985938 $Y=1949520
X1483 8612 8530 2 3 8585 AND2X1 $T=2209680 1803760 1 180 $X=2207040 $Y=1803358
X1484 424 5804 5808 2 5585 3 AOI2BB1X4 $T=1552980 1783600 0 0 $X=1552978 $Y=1783198
X1485 4394 220 2 219 114 4365 3 AOI22X1 $T=1254000 1793680 1 180 $X=1250700 $Y=1793278
X1486 4493 220 2 3789 68 4479 3 AOI22X1 $T=1277760 1793680 1 0 $X=1277758 $Y=1788240
X1487 5688 402 2 400 412 5685 3 AOI22X1 $T=1536480 1783600 0 180 $X=1533180 $Y=1778160
X1488 5772 5765 2 5743 5798 5800 3 AOI22X1 $T=1551000 1924720 0 0 $X=1550998 $Y=1924318
X1489 5951 5939 2 5900 5935 5902 3 AOI22X1 $T=1592580 1904560 1 180 $X=1589280 $Y=1904158
X1490 6379 487 2 488 489 6396 3 AOI22X1 $T=1694880 1985200 0 0 $X=1694878 $Y=1984798
X1491 514 487 2 488 450 6621 3 AOI22X1 $T=1752960 1975120 0 180 $X=1749660 $Y=1969680
X1492 490 528 2 527 559 573 3 AOI22X1 $T=1801800 1783600 0 0 $X=1801798 $Y=1783198
X1493 2383 101 2451 2455 3 2 2465 OAI2BB2X1 $T=826320 1965040 1 0 $X=826318 $Y=1959600
X1494 2636 113 2666 2663 3 2 2526 OAI2BB2X1 $T=877800 1834000 1 180 $X=873180 $Y=1833598
X1495 2818 68 2858 2859 3 2 2695 OAI2BB2X1 $T=917400 1934800 1 0 $X=917398 $Y=1929360
X1496 5975 319 5988 5986 3 2 5964 OAI2BB2X1 $T=1603140 1934800 1 180 $X=1598520 $Y=1934398
X1497 483 482 482 454 3 2 6237 OAI2BB2X1 $T=1683660 1813840 0 180 $X=1679040 $Y=1808400
X1498 485 482 482 419 3 2 6325 OAI2BB2X1 $T=1685640 1854160 1 180 $X=1681020 $Y=1853758
X1499 481 482 482 484 3 2 6398 OAI2BB2X1 $T=1683660 1864240 0 0 $X=1683658 $Y=1863838
X1500 825 738 10119 824 3 2 10099 OAI2BB2X1 $T=2541000 1985200 1 180 $X=2536380 $Y=1984798
X1501 3972 3969 3 2 221 XNOR2XL $T=1176120 1854160 1 180 $X=1170840 $Y=1853758
X1502 4261 4260 3 2 4235 XNOR2XL $T=1230900 1844080 1 180 $X=1225620 $Y=1843678
X1503 257 4307 3 2 4117 XNOR2XL $T=1241460 1965040 1 180 $X=1236180 $Y=1964638
X1504 4440 4439 3 2 3942 XNOR2XL $T=1266540 1864240 0 180 $X=1261260 $Y=1858800
X1505 6152 6221 3 2 471 XNOR2XL $T=1657260 1914640 1 180 $X=1651980 $Y=1914238
X1506 6292 6295 3 2 480 XNOR2XL $T=1673100 1934800 1 0 $X=1673098 $Y=1929360
X1507 7421 7422 3 2 6451 XNOR2XL $T=1941060 1975120 1 180 $X=1935780 $Y=1974718
X1508 8038 8055 3 2 666 XNOR2XL $T=2080980 1803760 0 180 $X=2075700 $Y=1798320
X1509 8090 8089 3 2 8055 XNOR2XL $T=2091540 1803760 0 180 $X=2086260 $Y=1798320
X1510 8364 700 3 2 8391 XNOR2XL $T=2148960 1813840 0 0 $X=2148958 $Y=1813438
X1511 8444 8443 3 2 688 XNOR2XL $T=2170080 1834000 1 180 $X=2164800 $Y=1833598
X1512 9376 9377 3 2 8920 XNOR2XL $T=2392500 1854160 1 180 $X=2387220 $Y=1853758
X1513 2498 118 2874 2 3 OR2X4 $T=920700 1803760 0 0 $X=920698 $Y=1803358
X1514 2317 121 2917 2 3 OR2X4 $T=943140 1793680 0 180 $X=939180 $Y=1788240
X1515 2840 133 3061 2 3 OR2X4 $T=964920 1844080 0 0 $X=964918 $Y=1843678
X1516 3414 3413 3357 2 3 OR2X4 $T=1052700 1823920 0 180 $X=1048740 $Y=1818480
X1517 3623 201 200 2 3 OR2X4 $T=1102200 1975120 0 180 $X=1098240 $Y=1969680
X1518 3056 4668 4615 2 3 OR2X4 $T=1319340 1813840 1 180 $X=1315380 $Y=1813438
X1519 577 576 6882 2 3 OR2X4 $T=1821600 1975120 0 180 $X=1817640 $Y=1969680
X1520 758 9167 8999 2 3 OR2X4 $T=2344980 1803760 0 180 $X=2341020 $Y=1798320
X1521 9492 9477 9456 2 3 OR2X4 $T=2410320 1904560 1 180 $X=2406360 $Y=1904158
X1522 9576 9274 9593 2 3 OR2X4 $T=2434740 1904560 1 0 $X=2434738 $Y=1899120
X1523 5216 350 5025 3 2 5086 OAI2BB1X4 $T=1435500 1783600 1 0 $X=1435498 $Y=1778160
X1524 365 333 5357 3 2 5271 OAI2BB1X4 $T=1462560 1783600 0 180 $X=1455960 $Y=1778160
X1525 791 9973 9974 3 2 10056 OAI2BB1X4 $T=2513280 1985200 1 0 $X=2513278 $Y=1979760
X1526 9977 10090 10087 3 2 10082 OAI2BB1X4 $T=2535720 1844080 1 180 $X=2529120 $Y=1843678
X1527 5453 385 3 2 INVX8 $T=1487640 1894480 1 0 $X=1487638 $Y=1889040
X1528 5557 397 3 2 INVX8 $T=1500180 1844080 0 0 $X=1500178 $Y=1843678
X1529 7316 618 3 2 INVX8 $T=1914660 1823920 0 180 $X=1910700 $Y=1818480
X1530 530 6751 3 2 INVX8 $T=2134440 1894480 1 0 $X=2134438 $Y=1889040
X1531 8980 747 3 2 INVX8 $T=2302740 1914640 0 180 $X=2298780 $Y=1909200
X1532 2197 2214 2213 3 2 NAND2BX2 $T=775500 1954960 0 180 $X=771540 $Y=1949520
X1533 9279 9325 9333 3 2 NAND2BX2 $T=2377980 1803760 0 0 $X=2377978 $Y=1803358
X1534 9634 9627 9527 3 2 NAND2BX2 $T=2443320 1954960 0 180 $X=2439360 $Y=1949520
X1535 160 3357 3432 3434 2 3 OAI2BB1X2 $T=1056000 1944880 1 0 $X=1055998 $Y=1939440
X1536 3458 174 155 3432 2 3 OAI2BB1X2 $T=1063920 1944880 1 0 $X=1063918 $Y=1939440
X1537 3521 190 3542 3546 2 3 OAI2BB1X2 $T=1081080 1874320 0 0 $X=1081078 $Y=1873918
X1538 3712 205 208 3716 2 3 OAI2BB1X2 $T=1117380 1965040 0 0 $X=1117378 $Y=1964638
X1539 461 149 6119 6139 2 3 OAI2BB1X2 $T=1634160 1793680 1 0 $X=1634158 $Y=1788240
X1540 8089 8038 8090 8129 2 3 OAI2BB1X2 $T=2094840 1793680 0 0 $X=2094838 $Y=1793278
X1541 690 8205 8214 8281 2 3 OAI2BB1X2 $T=2127180 1803760 1 0 $X=2127178 $Y=1798320
X1542 8364 8393 700 8429 2 3 OAI2BB1X2 $T=2157540 1813840 1 0 $X=2157538 $Y=1808400
X1543 9363 771 8622 9348 2 3 OAI2BB1X2 $T=2387220 1813840 0 180 $X=2382600 $Y=1808400
X1544 10064 10083 9976 10087 2 3 OAI2BB1X2 $T=2531100 1854160 0 0 $X=2531098 $Y=1853758
X1545 3658 3574 202 3 2 3623 AND3X2 $T=1103520 1975120 1 180 $X=1100220 $Y=1974718
X1546 4238 3813 4255 3 2 253 AND3X2 $T=1226940 1783600 1 0 $X=1226938 $Y=1778160
X1547 4283 4267 4281 3 2 255 AND3X2 $T=1234200 1793680 0 0 $X=1234198 $Y=1793278
X1548 4438 4430 4437 3 2 268 AND3X2 $T=1263900 1793680 0 0 $X=1263898 $Y=1793278
X1549 842 10082 10339 3 2 848 AND3X2 $T=2593140 1803760 1 0 $X=2593138 $Y=1798320
X1550 1970 71 2063 3 2 NOR2BX2 $T=728640 1954960 1 0 $X=728638 $Y=1949520
X1551 2947 3022 3 2 3103 XOR2XL $T=953700 1914640 0 0 $X=953698 $Y=1914238
X1552 185 176 3 2 3494 XOR2XL $T=1077780 1803760 1 180 $X=1072500 $Y=1803358
X1553 3807 3801 3 2 212 XOR2XL $T=1144440 1854160 1 180 $X=1139160 $Y=1853758
X1554 4045 4034 3 2 4025 XOR2XL $T=1191960 1904560 0 180 $X=1186680 $Y=1899120
X1555 4124 4144 3 2 4069 XOR2XL $T=1209120 1854160 1 180 $X=1203840 $Y=1853758
X1556 4366 4332 3 2 4394 XOR2XL $T=1249380 1844080 0 0 $X=1249378 $Y=1843678
X1557 4520 4519 3 2 4277 XOR2XL $T=1286340 1854160 1 180 $X=1281060 $Y=1853758
X1558 4632 4633 3 2 4410 XOR2XL $T=1310100 1834000 0 180 $X=1304820 $Y=1828560
X1559 6399 6400 3 2 6379 XOR2XL $T=1699500 1934800 0 180 $X=1694220 $Y=1929360
X1560 606 7235 3 2 6333 XOR2XL $T=1890240 1965040 0 180 $X=1884960 $Y=1959600
X1561 7367 7439 3 2 7416 XOR2XL $T=1942380 1864240 0 180 $X=1937100 $Y=1858800
X1562 7838 639 3 2 633 XOR2XL $T=2028840 1834000 1 180 $X=2023560 $Y=1833598
X1563 7998 7996 3 2 662 XOR2XL $T=2063160 1844080 0 180 $X=2057880 $Y=1838640
X1564 2 5082 4906 5086 5105 3 NAND3X2 $T=1405800 1793680 0 180 $X=1401180 $Y=1788240
X1565 2 5836 5809 5835 5671 3 NAND3X2 $T=1558920 1793680 1 0 $X=1558918 $Y=1788240
X1566 2 6066 6065 458 6061 3 NAND3X2 $T=1618320 1783600 0 0 $X=1618318 $Y=1783198
X1567 2 9624 9786 9794 9762 3 NAND3X2 $T=2473680 1864240 0 0 $X=2473678 $Y=1863838
X1568 122 123 125 3009 130 2 3 3044 SDFFRHQXL $T=946440 1954960 1 0 $X=946438 $Y=1949520
X1569 122 129 141 3101 130 2 3 3057 SDFFRHQXL $T=988020 1823920 0 180 $X=971520 $Y=1818480
X1570 122 123 128 3120 130 2 3 3084 SDFFRHQXL $T=988020 1954960 1 180 $X=971520 $Y=1954558
X1571 122 123 134 3123 130 2 3 3087 SDFFRHQXL $T=989340 1975120 0 180 $X=972840 $Y=1969680
X1572 122 123 146 3170 130 2 3 3244 SDFFRHQXL $T=995280 1954960 0 0 $X=995278 $Y=1954558
X1573 122 123 165 3331 130 2 3 3280 SDFFRHQXL $T=1049400 1965040 0 180 $X=1032900 $Y=1959600
X1574 122 123 155 224 216 2 3 3771 SDFFRHQXL $T=1187340 1985200 0 180 $X=1170840 $Y=1979760
X1575 122 123 190 4057 226 2 3 225 SDFFRHQXL $T=1202520 1965040 0 180 $X=1186020 $Y=1959600
X1576 122 129 4029 4118 226 2 3 227 SDFFRHQXL $T=1208460 1793680 1 180 $X=1191960 $Y=1793278
X1577 122 123 168 4232 226 2 3 4155 SDFFRHQXL $T=1229580 1965040 0 180 $X=1213080 $Y=1959600
X1578 277 123 271 270 226 2 3 4391 SDFFRHQXL $T=1278420 1965040 0 180 $X=1261920 $Y=1959600
X1579 277 123 302 4753 226 2 3 4844 SDFFRHQXL $T=1335840 1914640 0 0 $X=1335838 $Y=1914238
X1580 277 123 4863 4878 226 2 3 4843 SDFFRHQXL $T=1368840 1874320 0 180 $X=1352340 $Y=1868880
X1581 277 129 111 4906 226 2 3 4863 SDFFRHQXL $T=1372140 1793680 0 180 $X=1355640 $Y=1788240
X1582 277 123 372 5396 226 2 3 5261 SDFFRHQXL $T=1475100 1864240 1 180 $X=1458600 $Y=1863838
X1583 277 463 149 6044 226 2 3 6059 SDFFRHQXL $T=1638120 1834000 1 180 $X=1621620 $Y=1833598
X1584 277 465 462 6116 226 2 3 6078 SDFFRHQXL $T=1639440 1864240 1 180 $X=1622940 $Y=1863838
X1585 277 463 455 6139 226 2 3 6098 SDFFRHQXL $T=1644720 1823920 1 180 $X=1628220 $Y=1823518
X1586 277 465 470 6168 226 2 3 6134 SDFFRHQXL $T=1655280 1874320 0 180 $X=1638780 $Y=1868880
X1587 277 463 159 6237 226 2 3 6318 SDFFRHQXL $T=1655940 1813840 0 0 $X=1655938 $Y=1813438
X1588 277 463 148 476 226 2 3 6235 SDFFRHQXL $T=1675080 1803760 0 180 $X=1658580 $Y=1798320
X1589 277 465 481 6316 226 2 3 6261 SDFFRHQXL $T=1682340 1874320 1 180 $X=1665840 $Y=1873918
X1590 277 465 490 6325 226 2 3 6481 SDFFRHQXL $T=1694220 1854160 0 0 $X=1694218 $Y=1853758
X1591 277 465 485 6398 226 2 3 6467 SDFFRHQXL $T=1694220 1874320 0 0 $X=1694218 $Y=1873918
X1592 277 463 483 6444 226 2 3 496 SDFFRHQXL $T=1697520 1834000 0 0 $X=1697518 $Y=1833598
X1593 475 463 495 6065 226 2 3 6348 SDFFRHQXL $T=1714680 1793680 0 180 $X=1698180 $Y=1788240
X1594 277 465 500 6544 226 2 3 6580 SDFFRHQXL $T=1725240 1874320 0 0 $X=1725238 $Y=1873918
X1595 277 463 501 6556 226 2 3 509 SDFFRHQXL $T=1727880 1823920 0 0 $X=1727878 $Y=1823518
X1596 277 463 496 6557 226 2 3 501 SDFFRHQXL $T=1727880 1834000 0 0 $X=1727878 $Y=1833598
X1597 475 463 509 6601 504 2 3 503 SDFFRHQXL $T=1749660 1793680 0 180 $X=1733160 $Y=1788240
X1598 277 465 512 6597 226 2 3 520 SDFFRHQXL $T=1745700 1894480 0 0 $X=1745698 $Y=1894078
X1599 277 465 520 6673 226 2 3 500 SDFFRHQXL $T=1762200 1884400 1 180 $X=1745700 $Y=1883998
X1600 277 465 521 6675 226 2 3 6617 SDFFRHQXL $T=1763520 1914640 1 180 $X=1747020 $Y=1914238
X1601 475 463 523 6704 504 2 3 512 SDFFRHQXL $T=1769460 1783600 1 180 $X=1752960 $Y=1783198
X1602 277 465 530 6739 226 2 3 6779 SDFFRHQXL $T=1772760 1894480 0 0 $X=1772758 $Y=1894078
X1603 277 465 6753 6752 226 2 3 6788 SDFFRHQXL $T=1776060 1904560 0 0 $X=1776058 $Y=1904158
X1604 277 465 532 6891 226 2 3 6860 SDFFRHQXL $T=1818960 1894480 1 180 $X=1802460 $Y=1894078
X1605 277 465 574 6890 226 2 3 6878 SDFFRHQXL $T=1822260 1904560 1 180 $X=1805760 $Y=1904158
X1606 277 465 585 7004 226 2 3 574 SDFFRHQXL $T=1844700 1924720 1 180 $X=1828200 $Y=1924318
X1607 277 465 557 6941 226 2 3 7043 SDFFRHQXL $T=1830840 1894480 0 0 $X=1830838 $Y=1894078
X1608 277 465 575 7009 226 2 3 7119 SDFFRHQXL $T=1835460 1914640 0 0 $X=1835458 $Y=1914238
X1609 277 465 606 7204 226 2 3 597 SDFFRHQXL $T=1881000 1944880 1 180 $X=1864500 $Y=1944478
X1610 277 465 559 7207 226 2 3 7247 SDFFRHQXL $T=1879680 1904560 0 0 $X=1879678 $Y=1904158
X1611 277 465 597 7221 226 2 3 7249 SDFFRHQXL $T=1880340 1894480 0 0 $X=1880338 $Y=1894078
X1612 277 465 603 7187 226 2 3 7250 SDFFRHQXL $T=1880340 1934800 1 0 $X=1880338 $Y=1929360
X1613 277 465 613 7012 504 2 3 7261 SDFFRHQXL $T=1882980 1793680 0 0 $X=1882978 $Y=1793278
X1614 277 465 473 621 504 2 3 7541 SDFFRHQXL $T=1937100 1793680 0 0 $X=1937098 $Y=1793278
X1615 3044 2 128 3 BUFX3 $T=957660 1944880 1 180 $X=955020 $Y=1944478
X1616 123 2 129 3 BUFX3 $T=957660 1844080 0 0 $X=957658 $Y=1843678
X1617 3057 2 131 3 BUFX3 $T=965580 1823920 1 180 $X=962940 $Y=1823518
X1618 3084 2 134 3 BUFX3 $T=970200 1965040 1 0 $X=970198 $Y=1959600
X1619 3087 2 137 3 BUFX3 $T=975480 1975120 0 0 $X=975478 $Y=1974718
X1620 3244 2 141 3 BUFX3 $T=999240 1944880 1 180 $X=996600 $Y=1944478
X1621 3280 2 146 3 BUFX3 $T=1025640 1965040 0 180 $X=1023000 $Y=1959600
X1622 155 2 157 3 BUFX3 $T=1031580 1823920 0 0 $X=1031578 $Y=1823518
X1623 3771 2 165 3 BUFX3 $T=1134540 1985200 1 180 $X=1131900 $Y=1984798
X1624 130 2 216 3 BUFX3 $T=1141800 1944880 0 0 $X=1141798 $Y=1944478
X1625 205 2 248 3 BUFX3 $T=1224300 1813840 0 0 $X=1224298 $Y=1813438
X1626 4391 2 168 3 BUFX3 $T=1252680 1965040 0 180 $X=1250040 $Y=1959600
X1627 284 2 291 3 BUFX3 $T=1304820 1894480 0 0 $X=1304818 $Y=1894078
X1628 188 2 271 3 BUFX3 $T=1323300 1944880 0 0 $X=1323298 $Y=1944478
X1629 4843 2 302 3 BUFX3 $T=1354980 1904560 1 180 $X=1352340 $Y=1904158
X1630 329 2 333 3 BUFX3 $T=1397880 1783600 1 0 $X=1397878 $Y=1778160
X1631 5261 2 355 3 BUFX3 $T=1446720 1864240 1 180 $X=1444080 $Y=1863838
X1632 6059 2 372 3 BUFX3 $T=1617660 1834000 1 180 $X=1615020 $Y=1833598
X1633 6078 2 455 3 BUFX3 $T=1625580 1874320 1 0 $X=1625578 $Y=1868880
X1634 6098 2 149 3 BUFX3 $T=1634820 1823920 1 0 $X=1634818 $Y=1818480
X1635 6134 2 462 3 BUFX3 $T=1648020 1884400 1 0 $X=1648018 $Y=1878960
X1636 6235 2 159 3 BUFX3 $T=1658580 1793680 1 180 $X=1655940 $Y=1793278
X1637 6261 2 470 3 BUFX3 $T=1666500 1884400 1 0 $X=1666498 $Y=1878960
X1638 6318 2 483 3 BUFX3 $T=1679700 1823920 1 0 $X=1679698 $Y=1818480
X1639 6348 2 148 3 BUFX3 $T=1686960 1793680 0 180 $X=1684320 $Y=1788240
X1640 6467 2 481 3 BUFX3 $T=1705440 1884400 0 180 $X=1702800 $Y=1878960
X1641 6481 2 485 3 BUFX3 $T=1718640 1854160 0 0 $X=1718638 $Y=1853758
X1642 6580 2 490 3 BUFX3 $T=1731840 1854160 1 180 $X=1729200 $Y=1853758
X1643 6617 2 530 3 BUFX3 $T=1764180 1924720 0 0 $X=1764178 $Y=1924318
X1644 6860 2 557 3 BUFX3 $T=1801140 1894480 1 0 $X=1801138 $Y=1889040
X1645 6878 2 521 3 BUFX3 $T=1809720 1914640 0 0 $X=1809718 $Y=1914238
X1646 7220 2 7222 3 BUFX3 $T=1881660 1834000 0 0 $X=1881658 $Y=1833598
X1647 7250 2 596 3 BUFX3 $T=1888920 1924720 0 180 $X=1886280 $Y=1919280
X1648 7261 2 619 3 BUFX3 $T=1893540 1803760 0 180 $X=1890900 $Y=1798320
X1649 7249 2 611 3 BUFX3 $T=1896180 1874320 1 180 $X=1893540 $Y=1873918
X1650 7247 2 603 3 BUFX3 $T=1894200 1914640 0 0 $X=1894198 $Y=1914238
X1651 7541 2 7547 3 BUFX3 $T=1963500 1783600 0 0 $X=1963498 $Y=1783198
X1652 676 2 692 3 BUFX3 $T=2126520 1793680 1 0 $X=2126518 $Y=1788240
X1653 613 2 717 3 BUFX3 $T=2203740 1874320 0 180 $X=2201100 $Y=1868880
X1654 727 2 728 3 BUFX3 $T=2228160 1813840 1 0 $X=2228158 $Y=1808400
X1655 10412 10405 10405 2 10409 3 10431 10433 AOI221X1 $T=2611620 1793680 0 180 $X=2607000 $Y=1788240
X1656 6753 6798 6800 2 521 6789 3 6815 AOI32XL $T=1792560 1813840 0 0 $X=1792558 $Y=1813438
X1657 5720 406 2 3 CLKINVX4 $T=1521960 1793680 1 180 $X=1519320 $Y=1793278
X1658 5809 427 2 3 CLKINVX4 $T=1556280 1793680 1 0 $X=1556278 $Y=1788240
X1659 7032 582 2 3 CLKINVX4 $T=1848660 1854160 0 0 $X=1848658 $Y=1853758
X1660 7547 626 2 3 CLKINVX4 $T=1970100 1783600 1 0 $X=1970098 $Y=1778160
X1661 527 575 2 496 528 526 579 6465 3 AOI222X2 $T=1816980 1834000 0 0 $X=1816978 $Y=1833598
X1662 526 591 2 574 528 7024 582 7003 3 AOI222X2 $T=1851300 1834000 1 180 $X=1842060 $Y=1833598
X1663 606 527 2 596 528 614 526 7189 3 AOI222X2 $T=1882320 1844080 0 0 $X=1882318 $Y=1843678
X1664 210 2 112 3790 3 NOR2BXL $T=1123980 1793680 0 0 $X=1123978 $Y=1793278
X1665 426 2 5796 5748 3 NOR2BXL $T=1553640 1793680 1 180 $X=1551000 $Y=1793278
X1666 10227 2 10229 10271 3 NOR2BXL $T=2567400 1803760 0 0 $X=2567398 $Y=1803358
X1667 572 2 6862 6920 3 6942 NOR3BX1 $T=1816320 1803760 0 0 $X=1816318 $Y=1803358
X1668 7960 2 7926 7978 3 8001 NOR3BX1 $T=2061180 1783600 0 0 $X=2061178 $Y=1783198
X1669 7123 2 7121 6960 3 7048 7102 AOI211X1 $T=1857900 1844080 1 180 $X=1854600 $Y=1843678
X1670 7102 6982 7002 3 6942 7002 2 581 OAI32X1 $T=1842720 1803760 1 180 $X=1838100 $Y=1803358
X1671 7211 596 607 3 597 7234 2 7097 OAI32X1 $T=1885620 1864240 0 0 $X=1885618 $Y=1863838
X1672 2025 1997 3 2 2138 2135 AOI2BB1X1 $T=753060 1803760 1 0 $X=753058 $Y=1798320
X1673 2660 2731 3 2 2807 2823 AOI2BB1X1 $T=904200 1904560 1 0 $X=904198 $Y=1899120
X1674 5368 5321 3 2 5399 5473 AOI2BB1X1 $T=1472460 1934800 0 0 $X=1472458 $Y=1934398
X1675 8308 642 3 2 8272 8214 AOI2BB1X1 $T=2131140 1783600 0 180 $X=2127840 $Y=1778160
X1676 10229 10269 3 2 10266 847 AOI2BB1X1 $T=2568720 1793680 0 0 $X=2568718 $Y=1793278
X1677 3789 50 2 219 108 3942 3958 220 3 AOI222X1 $T=1164900 1783600 0 0 $X=1164898 $Y=1783198
X1678 527 532 2 528 501 6723 6559 526 3 AOI222X1 $T=1775400 1834000 1 180 $X=1770120 $Y=1833598
X1679 537 526 2 528 512 530 6697 527 3 AOI222X1 $T=1778040 1793680 0 180 $X=1772760 $Y=1788240
X1680 6753 527 2 528 503 533 6674 526 3 AOI222X1 $T=1778700 1803760 1 180 $X=1773420 $Y=1803358
X1681 526 612 2 597 528 527 7220 611 3 AOI222X1 $T=1884300 1834000 0 0 $X=1884298 $Y=1833598
X1682 3438 3450 172 3476 3 2 MXI2X1 $T=1058640 1975120 0 0 $X=1058638 $Y=1974718
X1683 3465 3494 183 3533 3 2 MXI2X1 $T=1069200 1793680 0 0 $X=1069198 $Y=1793278
X1684 8496 708 3 8530 2 8444 8525 OAI211X1 $T=2196480 1813840 1 180 $X=2192520 $Y=1813438
X1685 9494 9629 3 9609 2 9571 9615 OAI211X1 $T=2441340 1864240 1 180 $X=2437380 $Y=1863838
X1686 64 67 1965 3 2 1970 XNOR3X2 $T=708180 1965040 1 0 $X=708178 $Y=1959600
X1687 2614 2499 2634 3 2 2698 XNOR3X2 $T=862620 1944880 0 0 $X=862618 $Y=1944478
X1688 2663 2636 113 3 2 2592 XNOR3X2 $T=879780 1844080 0 180 $X=867900 $Y=1838640
X1689 2818 68 2859 3 2 2891 XNOR3X2 $T=915420 1924720 1 0 $X=915418 $Y=1919280
X1690 5986 5975 319 3 2 445 XNOR3X2 $T=1606440 1934800 0 180 $X=1594560 $Y=1929360
X1691 690 8214 8205 3 2 668 XNOR3X2 $T=2119920 1803760 1 180 $X=2108040 $Y=1803358
X1692 7547 692 8445 3 2 8393 XNOR3X2 $T=2160180 1793680 0 0 $X=2160178 $Y=1793278
X1693 772 775 776 3 2 9484 XNOR3X2 $T=2395800 1783600 1 0 $X=2395798 $Y=1778160
X1694 9706 9543 786 3 2 9538 XNOR3X2 $T=2450580 1844080 0 180 $X=2438700 $Y=1838640
X1695 804 810 812 3 2 9836 XNOR3X2 $T=2505360 1823920 0 0 $X=2505358 $Y=1823518
X1696 10083 9976 9977 3 2 9625 XNOR3X2 $T=2525820 1864240 0 180 $X=2513940 $Y=1858800
X1697 817 820 823 3 2 10083 XNOR3X2 $T=2527800 1803760 0 0 $X=2527798 $Y=1803358
X1698 840 839 10304 3 2 9472 XNOR3X2 $T=2591160 1793680 0 180 $X=2579280 $Y=1788240
X1699 50 2 3795 3795 150 3809 3 AOI22XL $T=1140480 1803760 1 0 $X=1140478 $Y=1798320
X1700 281 2 111 109 242 4177 3 AOI22XL $T=1266540 1783600 1 180 $X=1263240 $Y=1783198
X1701 5383 2 355 367 370 5387 3 AOI22XL $T=1465200 1823920 0 0 $X=1465198 $Y=1823518
X1702 5921 2 5932 5901 5974 5986 3 AOI22XL $T=1595880 1924720 1 0 $X=1595878 $Y=1919280
X1703 559 2 7206 603 7172 7121 3 AOI22XL $T=1871100 1844080 1 180 $X=1867800 $Y=1843678
X1704 185 192 3 3534 2 3533 AOI2BB1XL $T=1083720 1793680 1 180 $X=1080420 $Y=1793278
X1705 242 109 3 4177 2 3877 AOI2BB1XL $T=1214400 1783600 1 180 $X=1211100 $Y=1783198
X1706 7172 603 3 490 2 7206 AOI2BB1XL $T=1874400 1844080 1 0 $X=1874398 $Y=1838640
X1707 8527 8625 3 2 8525 8612 8622 OAI211X2 $T=2213640 1813840 1 180 $X=2207040 $Y=1813438
X1708 765 9348 3 2 9333 9356 9376 OAI211X2 $T=2381940 1803760 0 0 $X=2381938 $Y=1803358
X1709 9486 9538 3 2 9376 9504 9609 OAI211X2 $T=2423520 1844080 1 180 $X=2416920 $Y=1843678
X1710 9494 9629 3 2 9609 9571 9624 OAI211X2 $T=2442000 1864240 0 180 $X=2435400 $Y=1858800
X1711 8659 9027 9026 9019 2 3 739 AOI31X4 $T=2313960 1874320 1 180 $X=2308020 $Y=1873918
X1712 4844 180 3 2 BUFX4 $T=1347060 1914640 0 180 $X=1343760 $Y=1909200
X1713 321 233 3 2 BUFX4 $T=1370820 1904560 1 180 $X=1367520 $Y=1904158
X1714 382 5466 3 2 BUFX4 $T=1486980 1884400 1 0 $X=1486978 $Y=1878960
X1715 6788 532 3 2 BUFX4 $T=1790580 1914640 1 180 $X=1787280 $Y=1914238
X1716 594 592 3 2 BUFX4 $T=1854600 1985200 0 180 $X=1851300 $Y=1979760
X1717 6810 6806 550 2 6787 530 3 6861 AOI32X1 $T=1796520 1793680 1 0 $X=1796518 $Y=1788240
X1718 6893 6892 557 2 6863 532 3 6922 AOI32X1 $T=1812360 1844080 0 0 $X=1812358 $Y=1843678
X1719 575 7014 7008 2 582 6999 3 6961 AOI32X1 $T=1841400 1844080 1 180 $X=1836780 $Y=1843678
X1720 5692 5715 5568 3 5721 2 5766 OAI31X1 $T=1538460 1914640 1 0 $X=1538458 $Y=1909200
X1721 5837 5802 5568 3 5861 2 5875 OAI31X1 $T=1566840 1874320 0 0 $X=1566838 $Y=1873918
X1722 5846 5802 5568 3 5917 2 5931 OAI31X1 $T=1582020 1894480 0 0 $X=1582018 $Y=1894078
X1723 9138 9221 9114 3 9135 2 9273 OAI31X1 $T=2355540 1884400 1 0 $X=2355538 $Y=1878960
X1724 3452 3435 3436 3414 3 2 AND3X4 $T=1060620 1823920 0 180 $X=1056660 $Y=1818480
X1725 8445 7547 692 3 8473 2 OAI2BB1XL $T=2178660 1793680 1 0 $X=2178658 $Y=1788240
X1726 4031 3 58 2 CLKINVX8 $T=1195260 1823920 0 0 $X=1195258 $Y=1823518
X1727 242 3 62 2 CLKINVX8 $T=1209780 1823920 1 180 $X=1205820 $Y=1823518
X1728 4924 3 236 2 CLKINVX8 $T=1362900 1894480 1 180 $X=1358940 $Y=1894078
X1729 386 3 390 2 CLKINVX8 $T=1491600 1844080 0 0 $X=1491598 $Y=1843678
X1730 423 3 424 2 CLKINVX8 $T=1557600 1783600 1 0 $X=1557598 $Y=1778160
X1731 518 515 354 488 6681 487 542 3 2 AOI222X4 $T=1757580 1975120 1 0 $X=1757578 $Y=1969680
X1732 9045 8979 2 3 752 NOR2BX4 $T=2316600 1985200 1 0 $X=2316598 $Y=1979760
X1733 10339 10302 2 3 10409 NOR2BX4 $T=2588520 1803760 0 0 $X=2588518 $Y=1803358
X1734 5720 5740 5741 2 3 5748 NAND3BX2 $T=1542420 1793680 0 0 $X=1542418 $Y=1793278
X1735 247 236 233 3 218 2 231 230 3935 OAI222XL $T=1200540 1985200 0 180 $X=1195260 $Y=1979760
X1736 238 236 233 3 171 2 232 230 4057 OAI222XL $T=1201200 1985200 1 180 $X=1195920 $Y=1984798
X1737 196 233 236 3 252 2 254 230 4232 OAI222XL $T=1230900 1985200 1 0 $X=1230898 $Y=1979760
X1738 292 233 236 3 303 2 305 230 4651 OAI222XL $T=1338480 1934800 1 0 $X=1338478 $Y=1929360
X1739 310 236 233 3 307 2 306 230 4616 OAI222XL $T=1346400 1965040 0 180 $X=1341120 $Y=1959600
X1740 187 233 236 3 308 2 309 230 4753 OAI222XL $T=1342440 1924720 0 0 $X=1342438 $Y=1924318
X1741 319 236 233 3 317 2 316 230 4878 OAI222XL $T=1363560 1924720 1 180 $X=1358280 $Y=1924318
X1742 541 538 536 3 529 2 241 534 6739 OAI222XL $T=1780680 1874320 1 180 $X=1775400 $Y=1873918
X1743 535 536 538 3 6751 2 539 534 6675 OAI222XL $T=1776720 1864240 0 0 $X=1776718 $Y=1863838
X1744 6811 538 536 3 531 2 547 534 6752 OAI222XL $T=1795200 1884400 0 180 $X=1789920 $Y=1878960
X1745 6923 538 536 3 562 2 561 534 6891 OAI222XL $T=1813020 1874320 1 180 $X=1807740 $Y=1873918
X1746 7098 538 536 3 568 2 565 534 6890 OAI222XL $T=1815660 1884400 0 180 $X=1810380 $Y=1878960
X1747 6983 538 536 3 580 2 578 534 6941 OAI222XL $T=1825560 1874320 0 180 $X=1820280 $Y=1868880
X1748 589 538 536 3 587 2 586 534 7012 OAI222XL $T=1844700 1783600 1 180 $X=1839420 $Y=1783198
X1749 590 536 538 3 7032 2 588 534 7009 OAI222XL $T=1848000 1864240 1 180 $X=1842720 $Y=1863838
X1750 7129 538 536 3 595 2 593 534 7118 OAI222XL $T=1857900 1783600 1 180 $X=1852620 $Y=1783198
X1751 7173 538 536 3 598 2 452 534 7150 OAI222XL $T=1869120 1884400 0 180 $X=1863840 $Y=1878960
X1752 607 538 536 3 604 2 254 534 7144 OAI222XL $T=1875060 1864240 1 180 $X=1869780 $Y=1863838
X1753 7234 538 536 3 609 2 608 534 7221 OAI222XL $T=1883640 1874320 1 180 $X=1878360 $Y=1873918
X1754 7305 538 536 3 610 2 456 534 7207 OAI222XL $T=1883640 1884400 0 180 $X=1878360 $Y=1878960
X1755 4477 4479 3 2 274 AND2X4 $T=1274460 1793680 1 0 $X=1274458 $Y=1788240
X1756 6621 513 3 2 524 AND2X4 $T=1748340 1975120 0 0 $X=1748338 $Y=1974718
X1757 9795 790 3 2 9778 AND2X4 $T=2476320 1985200 0 180 $X=2473020 $Y=1979760
X1758 9920 9872 3 2 9868 AND2X4 $T=2501400 1954960 0 180 $X=2498100 $Y=1949520
X1759 136 138 134 3 2 3120 MX2X1 $T=976140 1934800 0 0 $X=976138 $Y=1934398
X1760 136 139 128 3 2 3009 MX2X1 $T=981420 1874320 0 180 $X=976140 $Y=1868880
X1761 136 140 131 3 2 3101 MX2X1 $T=982740 1793680 1 180 $X=977460 $Y=1793278
X1762 136 148 141 3 2 3170 MX2X1 $T=1002540 1934800 0 180 $X=997260 $Y=1929360
X1763 136 149 137 3 2 3123 MX2X1 $T=1003860 1934800 1 180 $X=998580 $Y=1934398
X1764 136 159 146 3 2 3331 MX2X1 $T=1041480 1934800 1 180 $X=1036200 $Y=1934398
X1765 5967 333 372 3 2 6044 MX2X1 $T=1597860 1834000 1 0 $X=1597858 $Y=1828560
X1766 5967 363 455 3 2 6116 MX2X1 $T=1613040 1844080 0 0 $X=1613038 $Y=1843678
X1767 5967 358 462 3 2 6168 MX2X1 $T=1652640 1864240 0 180 $X=1647360 $Y=1858800
X1768 5967 408 470 3 2 6316 MX2X1 $T=1665180 1864240 0 0 $X=1665178 $Y=1863838
X1769 126 130 3 2 INVX12 $T=952380 1975120 1 0 $X=952378 $Y=1969680
X1770 209 2 3 3789 BUFX8 $T=1133880 1783600 0 0 $X=1133878 $Y=1783198
X1771 402 5611 2 400 5603 5570 3 AOI22X2 $T=1516680 1793680 0 180 $X=1510740 $Y=1788240
X1772 216 226 3 2 BUFX16 $T=1176120 1944880 0 0 $X=1176118 $Y=1944478
X1773 4029 210 3 2 BUFX16 $T=1187340 1803760 0 0 $X=1187338 $Y=1803358
X1774 277 465 619 620 504 2 3 7368 SDFFRHQX1 $T=1910040 1793680 0 0 $X=1910038 $Y=1793278
X1775 277 465 7547 628 504 2 3 7569 SDFFRHQX1 $T=1962840 1793680 0 0 $X=1962838 $Y=1793278
X1776 3 2 292 ANTENNA $T=1337160 1934800 1 0 $X=1337158 $Y=1929360
X1777 277 123 284 4616 226 188 3 2 SDFFRHQX2 $T=1310100 1954960 0 180 $X=1290300 $Y=1949520
X1778 277 123 180 4651 226 284 3 2 SDFFRHQX2 $T=1317360 1934800 0 180 $X=1297560 $Y=1929360
X1779 3102 53 3 2 BUFX12 $T=979440 1783600 0 180 $X=972840 $Y=1778160
X1780 289 111 3 2 BUFX12 $T=1304820 1783600 1 0 $X=1304818 $Y=1778160
X1781 5500 393 3 2 BUFX12 $T=1493580 1854160 1 0 $X=1493578 $Y=1848720
X1782 122 164 123 3935 216 2 3 155 SDFFRHQX4 $T=1162260 1975120 1 0 $X=1162258 $Y=1969680
X1783 277 611 465 7118 504 2 3 550 SDFFRHQX4 $T=1881000 1783600 0 0 $X=1880998 $Y=1783198
X1784 475 625 465 634 504 2 3 639 SDFFRHQX4 $T=1990560 1793680 1 0 $X=1990558 $Y=1788240
X1785 122 129 50 151 130 143 3102 3 2 SDFFRX4 $T=1010460 1783600 0 180 $X=987360 $Y=1778160
X1786 122 129 68 229 226 242 243 3 2 SDFFRX4 $T=1186680 1834000 0 0 $X=1186678 $Y=1833598
X1787 122 129 242 240 226 4031 4029 3 2 SDFFRX4 $T=1210440 1813840 0 180 $X=1187340 $Y=1808400
X1788 277 465 7119 7150 226 10479 559 3 2 SDFFRX4 $T=1860540 1914640 0 0 $X=1860538 $Y=1914238
X1789 277 465 596 7144 226 10480 606 3 2 SDFFRX4 $T=1861200 1944880 1 0 $X=1861198 $Y=1939440
X1790 527 2 3 7024 BUFX2 $T=1839420 1834000 0 0 $X=1839418 $Y=1833598
X1791 6143 3 463 2 CLKINVX2 $T=1642080 1834000 0 0 $X=1642078 $Y=1833598
X1792 6143 3 465 2 CLKINVX2 $T=1644720 1854160 0 0 $X=1644718 $Y=1853758
X1793 1841 50 68 2 3 57 CMPR22X1 $T=724680 1914640 0 180 $X=716760 $Y=1909200
X1794 8167 6983 7098 2 3 8188 CMPR22X1 $T=2096160 1924720 1 0 $X=2096158 $Y=1919280
X1795 2272 2197 3 85 2195 2205 2 AOI2BB2X2 $T=774180 1965040 1 180 $X=768240 $Y=1964638
X1796 616 610 3 610 616 7316 2 AOI2BB2X2 $T=1910700 1823920 0 180 $X=1904760 $Y=1818480
X1797 2818 53 58 2 3 2750 ADDHX1 $T=910800 1944880 0 180 $X=902880 $Y=1939440
X1798 278 3 2 122 CLKBUFX20 $T=1285020 1844080 0 180 $X=1269180 $Y=1838640
X1799 278 3 2 277 CLKBUFX20 $T=1277100 1954960 0 0 $X=1277098 $Y=1954558
X1800 278 3 2 475 CLKBUFX20 $T=1657260 1803760 0 0 $X=1657258 $Y=1803358
X1801 5322 354 356 353 5214 5199 346 3 2 5173 CMPR42X1 $T=1448040 1985200 0 180 $X=1425600 $Y=1979760
X1802 375 371 373 5234 362 5339 5322 3 2 5236 CMPR42X1 $T=1473120 1985200 1 180 $X=1450680 $Y=1984798
X1803 8112 7407 550 7032 6811 8211 8188 3 2 8212 CMPR42X1 $T=2095500 1924720 0 0 $X=2095498 $Y=1924318
X1804 8309 6923 541 7129 8326 8310 8112 3 2 8273 CMPR42X1 $T=2154900 1934800 0 180 $X=2132460 $Y=1929360
X1805 8392 6811 702 8338 8313 8315 8309 3 2 8288 CMPR42X1 $T=2156880 1904560 1 180 $X=2134440 $Y=1904158
X1806 8493 7129 589 8412 8411 8397 8392 3 2 8365 CMPR42X1 $T=2172720 1894480 0 180 $X=2150280 $Y=1889040
X1807 8487 7129 709 8474 8540 8582 8583 3 2 8541 CMPR42X1 $T=2182620 1924720 0 0 $X=2182618 $Y=1924318
X1808 8583 718 7098 8539 8537 8512 8493 3 2 8495 CMPR42X1 $T=2209020 1894480 0 180 $X=2186580 $Y=1889040
X1809 8781 589 719 8616 8469 8599 8487 3 2 8584 CMPR42X1 $T=2223540 1934800 1 180 $X=2201100 $Y=1934398
X1810 8695 702 729 8725 8710 8776 8703 3 2 8869 CMPR42X1 $T=2235420 1864240 0 0 $X=2235418 $Y=1863838
X1811 8696 702 718 8475 8743 8777 8781 3 2 8798 CMPR42X1 $T=2235420 1944880 1 0 $X=2235418 $Y=1939440
X1812 8703 719 6751 8726 8772 8778 8708 3 2 8889 CMPR42X1 $T=2236080 1884400 1 0 $X=2236078 $Y=1878960
X1813 8705 713 521 589 8773 8780 8695 3 2 8800 CMPR42X1 $T=2236740 1844080 0 0 $X=2236738 $Y=1843678
X1814 8708 7129 709 8672 8621 8783 8714 3 2 8833 CMPR42X1 $T=2237400 1894480 0 0 $X=2237398 $Y=1894078
X1815 8711 589 709 8676 8601 8795 8696 3 2 8814 CMPR42X1 $T=2238060 1924720 0 0 $X=2238058 $Y=1924318
X1816 8714 718 729 8598 8641 8797 8711 3 2 8832 CMPR42X1 $T=2238720 1904560 0 0 $X=2238718 $Y=1904158
X1817 9221 9114 3 9223 9174 9173 2 OAI31XL $T=2354880 1874320 0 180 $X=2350920 $Y=1868880
.ENDS
***************************************
.SUBCKT ICV_68 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
** N=68 EP=38 IP=96 FDC=0
X24 3 21 PDO12CDG $T=793200 0 0 0 $X=795518 $Y=598
X25 4 31 PDO12CDG $T=872975 0 0 0 $X=875293 $Y=598
X26 5 22 PDO12CDG $T=952750 0 0 0 $X=955068 $Y=598
X27 6 32 PDO12CDG $T=1032525 0 0 0 $X=1034843 $Y=598
X28 7 23 PDO12CDG $T=1112300 0 0 0 $X=1114618 $Y=598
X29 8 24 PDO12CDG $T=1271845 0 0 0 $X=1274163 $Y=598
X30 9 33 PDO12CDG $T=1351615 0 0 0 $X=1353933 $Y=598
X31 10 34 PDO12CDG $T=1511155 0 0 0 $X=1513473 $Y=598
X32 11 35 PDO12CDG $T=1670695 0 0 0 $X=1673013 $Y=598
X33 12 25 PDO12CDG $T=1750465 0 0 0 $X=1752783 $Y=598
X34 13 36 PDO12CDG $T=1830235 0 0 0 $X=1832553 $Y=598
X35 14 26 PDO12CDG $T=1910005 0 0 0 $X=1912323 $Y=598
X36 15 27 PDO12CDG $T=2069545 0 0 0 $X=2071863 $Y=598
X37 16 28 PDO12CDG $T=2229095 0 0 0 $X=2231413 $Y=598
X38 17 37 PDO12CDG $T=2308870 0 0 0 $X=2311188 $Y=598
X39 18 29 PDO12CDG $T=2388645 0 0 0 $X=2390963 $Y=598
X40 19 38 PDO12CDG $T=2468420 0 0 0 $X=2470738 $Y=598
X41 20 30 PDO12CDG $T=2548195 0 0 0 $X=2550513 $Y=598
.ENDS
***************************************
.SUBCKT ICV_67
** N=26959 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_66
** N=27820 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_65 2 4 88 90 91 93 95 103 104 106 107 108 110 113 115 117 119 121 122 124
+ 125 128 131 132 138 139 140 143 144 145 146 148 151 153 155 157 158 161 1421 1422
** N=23885 EP=40 IP=632 FDC=0
X0 110 4 3944 2 3946 NAND2X1 $T=1428900 735280 1 0 $X=1428898 $Y=729840
X1 3931 4 3976 2 3991 NAND2X1 $T=1438140 715120 0 0 $X=1438138 $Y=714718
X2 115 4 3993 2 4073 NAND2X1 $T=1455960 735280 0 180 $X=1453980 $Y=729840
X3 4080 4 121 2 4171 NAND2X1 $T=1492920 735280 1 0 $X=1492918 $Y=729840
X4 4011 4 4225 2 4317 NAND2X1 $T=1534500 705040 0 0 $X=1534498 $Y=704638
X5 131 4 4288 2 132 NAND2X1 $T=1535160 725200 0 0 $X=1535158 $Y=724798
X6 4318 4 4317 2 4319 NAND2X1 $T=1543740 705040 0 0 $X=1543738 $Y=704638
X7 3748 4 4319 2 4501 NAND2X1 $T=1568820 715120 0 0 $X=1568818 $Y=714718
X8 3733 4 4393 2 4439 NAND2X1 $T=1568820 735280 0 0 $X=1568818 $Y=734878
X9 145 4 153 2 4652 NAND2X1 $T=1647360 735280 0 0 $X=1647358 $Y=734878
X10 155 4 153 2 4713 NAND2X1 $T=1653960 735280 0 0 $X=1653958 $Y=734878
X11 3734 2 4 4206 138 NOR2X4 $T=1584000 725200 1 180 $X=1579380 $Y=724798
X12 4526 4 4501 4553 2 NAND2BX1 $T=1607760 725200 1 0 $X=1607758 $Y=719760
X13 138 4 140 4680 2 NAND2BX1 $T=1634160 725200 0 0 $X=1634158 $Y=724798
X14 132 4526 4 4501 2 4525 OAI21X1 $T=1603140 725200 1 180 $X=1599840 $Y=724798
X15 3929 4 3928 3873 2 3945 OAI21XL $T=1420980 715120 0 0 $X=1420978 $Y=714718
X16 4040 4 3991 3975 2 3995 OAI21XL $T=1448040 715120 1 180 $X=1445400 $Y=714718
X17 3930 4 4040 3928 2 4053 OAI21XL $T=1458600 715120 0 0 $X=1458598 $Y=714718
X18 4126 4 122 4070 2 4152 OAI21XL $T=1487640 725200 1 0 $X=1487638 $Y=719760
X19 4135 4 122 4052 2 4134 OAI21XL $T=1490280 705040 1 180 $X=1487640 $Y=704638
X20 4155 4 122 4108 2 4208 OAI21XL $T=1495560 715120 0 0 $X=1495558 $Y=714718
X21 4171 4 122 4081 2 4195 OAI21XL $T=1500180 735280 1 0 $X=1500178 $Y=729840
X22 140 4 4410 4439 2 4484 OAI21XL $T=1591920 735280 0 0 $X=1591918 $Y=734878
X23 3961 4 2 3960 INVX1 $T=1434840 725200 0 180 $X=1433520 $Y=719760
X24 4041 4 2 4040 INVX1 $T=1451340 725200 1 0 $X=1451338 $Y=719760
X25 4073 4 2 4080 INVX1 $T=1463220 735280 1 0 $X=1463218 $Y=729840
X26 4227 4 2 4393 INVX1 $T=1564200 725200 1 0 $X=1564198 $Y=719760
X27 4439 4 2 4451 INVX1 $T=1579380 735280 0 0 $X=1579378 $Y=734878
X28 145 4 2 146 INVX1 $T=1607100 735280 0 180 $X=1605780 $Y=729840
X29 4525 4 2 148 INVX1 $T=1618980 735280 1 0 $X=1618978 $Y=729840
X30 2 107 3901 3930 4 NOR2X1 $T=1419660 725200 1 0 $X=1419658 $Y=719760
X31 2 3929 3930 3976 4 NOR2X1 $T=1431540 715120 1 0 $X=1431538 $Y=709680
X32 2 3930 4073 4071 4 NOR2X1 $T=1464540 705040 0 0 $X=1464538 $Y=704638
X33 2 4135 124 4154 4 NOR2X1 $T=1492920 705040 0 0 $X=1492918 $Y=704638
X34 2 4134 4211 4225 4 NOR2X1 $T=1510080 705040 0 0 $X=1510078 $Y=704638
X35 2 131 4288 4367 4 NOR2X1 $T=1535820 715120 0 0 $X=1535818 $Y=714718
X36 2 4410 138 143 4 NOR2X1 $T=1597860 735280 0 0 $X=1597858 $Y=734878
X37 4319 3748 4 2 4526 NOR2X2 $T=1556280 715120 0 0 $X=1556278 $Y=714718
X38 4393 3733 4 2 4410 NOR2X2 $T=1561560 735280 0 0 $X=1561558 $Y=734878
X39 4367 4526 4 2 145 NOR2X2 $T=1605120 715120 0 0 $X=1605118 $Y=714718
X40 108 103 4 2 3931 OR2XL $T=1422300 725200 1 0 $X=1422298 $Y=719760
X41 4206 3734 140 4 2 NAND2X2 $T=1593240 725200 1 180 $X=1589940 $Y=724798
X42 3931 2 3961 4 3994 AND2X2 $T=1440120 725200 1 0 $X=1440118 $Y=719760
X43 3944 110 4 2 3993 OR2X2 $T=1436160 735280 1 0 $X=1436158 $Y=729840
X44 4225 4011 4 2 4318 OR2X2 $T=1525260 705040 0 0 $X=1525258 $Y=704638
X45 4410 4451 4 2 139 OR2X2 $T=1586640 735280 0 0 $X=1586638 $Y=734878
X46 103 4 2 104 3873 NAND2XL $T=1401180 725200 0 0 $X=1401178 $Y=724798
X47 107 4 2 3901 3928 NAND2XL $T=1411740 725200 1 0 $X=1411738 $Y=719760
X48 103 4 2 108 3961 NAND2XL $T=1430220 725200 0 0 $X=1430218 $Y=724798
X49 3946 4 2 3993 4010 NAND2XL $T=1443420 735280 1 0 $X=1443418 $Y=729840
X50 4071 4 2 121 4135 NAND2XL $T=1479720 715120 1 0 $X=1479718 $Y=709680
X51 4072 4 2 121 4126 NAND2XL $T=1479720 715120 0 0 $X=1479718 $Y=714718
X52 4099 4 2 121 4155 NAND2XL $T=1485000 715120 0 0 $X=1484998 $Y=714718
X53 93 3733 4 2 INVX4 $T=1351680 735280 0 0 $X=1351678 $Y=734878
X54 4080 117 2 4041 4081 4 AOI21X1 $T=1469160 735280 0 180 $X=1466520 $Y=729840
X55 125 4228 2 4195 4241 4 AOI21X1 $T=1516020 735280 1 0 $X=1516018 $Y=729840
X56 4525 143 2 4484 144 4 AOI21X1 $T=1606440 735280 1 180 $X=1603800 $Y=734878
X57 145 151 2 4525 4592 4 AOI21X1 $T=1634160 735280 0 180 $X=1631520 $Y=729840
X58 155 151 2 4682 4681 4 AOI21X1 $T=1655280 725200 1 180 $X=1652640 $Y=724798
X59 157 4652 4 4592 2 4651 OAI21X2 $T=1649340 735280 0 180 $X=1644060 $Y=729840
X60 157 4713 4 4681 2 4714 OAI21X2 $T=1661880 735280 1 0 $X=1661878 $Y=729840
X61 4553 4714 158 4 2 XNOR2X4 $T=1661220 725200 1 0 $X=1661218 $Y=719760
X62 4680 4651 161 4 2 XNOR2X4 $T=1677060 725200 0 0 $X=1677058 $Y=724798
X63 95 4 3734 2 INVX2 $T=1354320 725200 0 0 $X=1354318 $Y=724798
X64 4367 4 155 2 INVX2 $T=1618320 715120 0 0 $X=1618318 $Y=714718
X65 132 2 4 4682 INVXL $T=1647360 725200 1 0 $X=1647358 $Y=719760
X66 4010 119 4 2 128 XOR2X1 $T=1475100 735280 0 0 $X=1475098 $Y=734878
X67 4009 4241 4 2 4288 XOR2X1 $T=1516020 725200 1 0 $X=1516018 $Y=719760
X68 3873 2 3929 4011 4 NOR2BX1 $T=1423620 705040 0 0 $X=1423618 $Y=704638
X69 3976 2 4073 4072 4 NOR2BX1 $T=1469160 725200 1 0 $X=1469158 $Y=719760
X70 103 106 108 3901 2 4 3944 ADDFX2 $T=1407120 735280 1 0 $X=1407118 $Y=729840
X71 3994 4170 4 2 4206 XNOR2X1 $T=1498200 725200 1 0 $X=1498198 $Y=719760
X72 2 103 104 3929 4 NOR2XL $T=1401180 715120 0 0 $X=1401178 $Y=714718
X73 2 4073 3991 4099 4 NOR2XL $T=1464540 715120 0 0 $X=1464538 $Y=714718
X74 2 4126 124 4153 4 NOR2XL $T=1490280 715120 0 0 $X=1490278 $Y=714718
X75 2 4171 124 4228 4 NOR2XL $T=1504140 735280 1 0 $X=1504138 $Y=729840
X76 2 4155 124 4207 4 NOR2XL $T=1506120 715120 1 0 $X=1506118 $Y=709680
X77 88 90 91 4 2 3589 XOR3X2 $T=1304820 715120 0 0 $X=1304818 $Y=714718
X78 3931 3945 2 3960 4 3975 AOI21XL $T=1429560 715120 0 0 $X=1429558 $Y=714718
X79 4071 117 2 4053 4 4052 AOI21XL $T=1461240 715120 0 180 $X=1458600 $Y=709680
X80 4099 117 2 3995 4 4108 AOI21XL $T=1471800 715120 0 0 $X=1471798 $Y=714718
X81 125 4153 2 4152 4 4170 AOI21XL $T=1492920 725200 1 0 $X=1492918 $Y=719760
X82 125 4207 2 4208 4 4227 AOI21XL $T=1506780 725200 1 0 $X=1506778 $Y=719760
X83 113 3993 3946 4 4041 2 OAI2BB1X1 $T=1448040 735280 1 0 $X=1448038 $Y=729840
X84 3930 4 3928 2 4009 NAND2BXL $T=1445400 725200 1 0 $X=1445398 $Y=719760
X85 3589 2 3748 4 CLKINVX3 $T=1338480 715120 0 0 $X=1338478 $Y=714718
X86 4154 125 2 4 4211 AND2X1 $T=1501500 705040 0 0 $X=1501498 $Y=704638
X87 3976 4041 117 2 4072 4 3945 4070 AOI221X1 $T=1466520 725200 0 180 $X=1461900 $Y=719760
.ENDS
***************************************
.SUBCKT AOI32X2 A0 A1 A2 VDD B1 B0 Y VSS
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND4X2 A B C D VSS VDD Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI31X4 B0 A0 A1 A2 Y VDD VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4X2 A B VDD D C VSS Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI32X4 B1 B0 A0 A1 A2 VDD Y VSS
** N=10 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_64 1 3 42 43 44 45 46 47 48 49 50 51 52 53 56 57 62 63 64 65
+ 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85
+ 86 87 89 91 93 95 96 97 99 100 102 103 104 108 109 110 111 112 113 114
+ 115 116 117 118 119 120 122 123 124 125 126 127 128 129 130 131 132 133 134 135
+ 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155
+ 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175
+ 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195
+ 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215
+ 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 236 237
+ 239 240 241 242 243 244 245 246 247 248 255 257 258 259 260 261 262 263 264 265
+ 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285
+ 342 343 344 345 346 347 348 349 350 351 1369 1370
** N=34202 EP=232 IP=7189 FDC=0
X0 2695 3 2615 1 2592 NAND2X1 $T=944460 916720 1 180 $X=942480 $Y=916318
X1 2799 3 2712 1 2734 NAND2X1 $T=973500 936880 1 180 $X=971520 $Y=936478
X2 2841 3 2825 1 2798 NAND2X1 $T=987360 916720 0 180 $X=985380 $Y=911280
X3 2884 3 2886 1 2735 NAND2X1 $T=1001220 946960 1 0 $X=1001218 $Y=941520
X4 3594 3 3428 1 3644 NAND2X1 $T=1163580 957040 1 0 $X=1163578 $Y=951600
X5 3361 3 3424 1 3791 NAND2X1 $T=1168860 836080 0 0 $X=1168858 $Y=835678
X6 3339 3 3691 1 3706 NAND2X1 $T=1176780 826000 1 0 $X=1176778 $Y=820560
X7 3711 3 3717 1 3743 NAND2X1 $T=1183380 785680 0 0 $X=1183378 $Y=785278
X8 3802 3 3847 1 4051 NAND2X1 $T=1211100 765520 1 0 $X=1211098 $Y=760080
X9 3849 3 3848 1 4076 NAND2X1 $T=1234200 765520 0 0 $X=1234198 $Y=765118
X10 4047 3 4091 1 4107 NAND2X1 $T=1241460 916720 0 0 $X=1241458 $Y=916318
X11 4080 3 109 1 4172 NAND2X1 $T=1250040 967120 0 0 $X=1250038 $Y=966718
X12 4414 3 4359 1 4436 NAND2X1 $T=1315380 755440 0 0 $X=1315378 $Y=755038
X13 144 3 134 1 140 NAND2X1 $T=1396560 977200 0 0 $X=1396558 $Y=976798
X14 141 3 134 1 4811 NAND2X1 $T=1397220 967120 0 0 $X=1397218 $Y=966718
X15 4944 3 4947 1 5022 NAND2X1 $T=1418340 826000 0 0 $X=1418338 $Y=825598
X16 4981 3 4921 1 4994 NAND2X1 $T=1426260 785680 0 0 $X=1426258 $Y=785278
X17 4984 3 4987 1 4993 NAND2X1 $T=1427580 745360 0 0 $X=1427578 $Y=744958
X18 4966 3 4923 1 5039 NAND2X1 $T=1432860 775600 0 0 $X=1432858 $Y=775198
X19 5023 3 4968 1 5029 NAND2X1 $T=1436820 836080 0 0 $X=1436818 $Y=835678
X20 5039 3 5053 1 5122 NAND2X1 $T=1443420 785680 0 0 $X=1443418 $Y=785278
X21 5006 3 5069 1 5139 NAND2X1 $T=1446060 775600 0 0 $X=1446058 $Y=775198
X22 5053 3 5136 1 5155 NAND2X1 $T=1456620 785680 0 0 $X=1456618 $Y=785278
X23 5055 3 5116 1 5161 NAND2X1 $T=1457940 856240 1 0 $X=1457938 $Y=850800
X24 5069 3 5053 1 5154 NAND2X1 $T=1459260 775600 0 0 $X=1459258 $Y=775198
X25 5175 3 5123 1 5176 NAND2X1 $T=1467180 876400 0 180 $X=1465200 $Y=870960
X26 148 3 153 1 5178 NAND2X1 $T=1469820 745360 0 0 $X=1469818 $Y=744958
X27 5008 3 5118 1 5302 NAND2X1 $T=1471140 967120 0 0 $X=1471138 $Y=966718
X28 5163 3 5220 1 5244 NAND2X1 $T=1479060 926800 0 180 $X=1477080 $Y=921360
X29 5176 3 5238 1 5286 NAND2X1 $T=1481040 886480 1 0 $X=1481038 $Y=881040
X30 5072 3 5282 1 5278 NAND2X1 $T=1490940 936880 1 0 $X=1490938 $Y=931440
X31 156 3 5203 1 157 NAND2X1 $T=1498200 977200 1 180 $X=1496220 $Y=976798
X32 153 3 5318 1 5365 NAND2X1 $T=1498200 765520 0 0 $X=1498198 $Y=765118
X33 5379 3 5326 1 5320 NAND2X1 $T=1500840 936880 1 180 $X=1498860 $Y=936478
X34 5314 3 5365 1 5297 NAND2X1 $T=1506120 765520 0 0 $X=1506118 $Y=765118
X35 4452 3 5400 1 5452 NAND2X1 $T=1516680 815920 0 0 $X=1516678 $Y=815518
X36 4439 3 5430 1 5523 NAND2X1 $T=1519320 846160 1 180 $X=1517340 $Y=845758
X37 4193 3 5429 1 5516 NAND2X1 $T=1519320 755440 0 0 $X=1519318 $Y=755038
X38 4494 3 162 1 5474 NAND2X1 $T=1527240 745360 0 0 $X=1527238 $Y=744958
X39 4715 3 5364 1 5498 NAND2X1 $T=1531200 826000 0 0 $X=1531198 $Y=825598
X40 4417 3 5402 1 5674 NAND2X1 $T=1554300 896560 1 180 $X=1552320 $Y=896158
X41 4312 3 5547 1 5680 NAND2X1 $T=1554300 926800 0 180 $X=1552320 $Y=921360
X42 4453 3 5627 1 5656 NAND2X1 $T=1554300 957040 1 0 $X=1554298 $Y=951600
X43 5717 3 5548 1 5713 NAND2X1 $T=1571460 967120 0 180 $X=1569480 $Y=961680
X44 5538 3 5675 1 5726 NAND2X1 $T=1572120 886480 0 0 $X=1572118 $Y=886078
X45 5498 3 5774 1 5759 NAND2X1 $T=1583340 846160 1 0 $X=1583338 $Y=840720
X46 5680 3 5760 1 5775 NAND2X1 $T=1584660 926800 1 0 $X=1584658 $Y=921360
X47 5758 3 5787 1 5845 NAND2X1 $T=1592580 765520 0 0 $X=1592578 $Y=765118
X48 5656 3 5717 1 5896 NAND2X1 $T=1595220 957040 1 0 $X=1595218 $Y=951600
X49 6069 3 192 1 6162 NAND2X1 $T=1657920 745360 0 0 $X=1657918 $Y=744958
X50 6901 3 5963 1 6900 NAND2X1 $T=1822920 926800 0 180 $X=1820940 $Y=921360
X51 7102 3 5964 1 7061 NAND2X1 $T=1857240 957040 0 180 $X=1855260 $Y=951600
X52 5962 3 7148 1 7192 NAND2X1 $T=1877700 856240 0 0 $X=1877698 $Y=855838
X53 7231 3 7213 1 7237 NAND2X1 $T=1892880 906640 1 180 $X=1890900 $Y=906238
X54 7233 3 7235 1 7257 NAND2X1 $T=1894860 896560 1 0 $X=1894858 $Y=891120
X55 7215 3 7177 1 227 NAND2X1 $T=1895520 967120 0 0 $X=1895518 $Y=966718
X56 5932 3 7234 1 7215 NAND2X1 $T=1899480 957040 0 0 $X=1899478 $Y=956638
X57 6193 3 7317 1 7298 NAND2X1 $T=1909380 815920 1 0 $X=1909378 $Y=810480
X58 7408 3 7427 1 7452 NAND2X1 $T=1945680 886480 0 0 $X=1945678 $Y=886078
X59 6167 3 7553 1 7533 NAND2X1 $T=1966140 795760 0 0 $X=1966138 $Y=795358
X60 6668 3 7667 1 7669 NAND2X1 $T=1981980 916720 0 0 $X=1981978 $Y=916318
X61 7669 3 7723 1 7714 NAND2X1 $T=1995180 926800 1 0 $X=1995178 $Y=921360
X62 7877 3 7875 1 7876 NAND2X1 $T=2020260 957040 1 0 $X=2020258 $Y=951600
X63 7897 3 7880 1 7895 NAND2X1 $T=2026200 846160 0 180 $X=2024220 $Y=840720
X64 7946 3 7880 1 7150 NAND2X1 $T=2040060 896560 0 0 $X=2040058 $Y=896158
X65 8122 3 8117 1 8113 NAND2X1 $T=2075700 906640 1 180 $X=2073720 $Y=906238
X66 8268 3 8305 1 8161 NAND2X1 $T=2110020 876400 0 0 $X=2110018 $Y=875998
X67 8385 3 8327 1 8200 NAND2X1 $T=2127840 846160 1 180 $X=2125860 $Y=845758
X68 8387 3 8393 1 8324 NAND2X1 $T=2131140 876400 0 0 $X=2131138 $Y=875998
X69 8445 3 8462 1 8385 NAND2X1 $T=2148960 876400 1 180 $X=2146980 $Y=875998
X70 8389 3 8443 1 8458 NAND2X1 $T=2149620 886480 0 0 $X=2149618 $Y=886078
X71 271 3 270 1 8545 NAND2X1 $T=2175360 977200 1 180 $X=2173380 $Y=976798
X72 8657 3 8632 1 8637 NAND2X1 $T=2185260 856240 1 180 $X=2183280 $Y=855838
X73 270 3 8499 1 342 NAND2X1 $T=2185920 977200 0 0 $X=2185918 $Y=976798
X74 8674 3 8657 1 8616 NAND2X1 $T=2193180 876400 0 180 $X=2191200 $Y=870960
X75 8766 3 8632 1 8764 NAND2X1 $T=2209020 856240 1 180 $X=2207040 $Y=855838
X76 278 3 8810 1 8745 NAND2X1 $T=2216280 967120 0 0 $X=2216278 $Y=966718
X77 8836 3 8829 1 8574 NAND2X1 $T=2222220 866320 0 180 $X=2220240 $Y=860880
X78 8851 3 8792 1 8746 NAND2X1 $T=2227500 886480 1 180 $X=2225520 $Y=886078
X79 8859 3 8914 1 8899 NAND2X1 $T=2242020 876400 0 180 $X=2240040 $Y=870960
X80 8860 3 8943 1 8836 NAND2X1 $T=2259180 876400 1 0 $X=2259178 $Y=870960
X81 5455 1 3 5513 5540 NOR2X4 $T=1544400 836080 1 180 $X=1539780 $Y=835678
X82 4416 1 3 5410 5672 NOR2X4 $T=1550340 775600 0 0 $X=1550338 $Y=775198
X83 5625 1 3 5521 5590 NOR2X4 $T=1554960 866320 0 180 $X=1550340 $Y=860880
X84 7388 1 3 7493 7526 NOR2X4 $T=1952280 795760 1 180 $X=1947660 $Y=795358
X85 6167 1 3 7553 7493 NOR2X4 $T=1956240 795760 1 0 $X=1956238 $Y=790320
X86 6273 1 3 7637 7598 NOR2X4 $T=1976700 886480 1 0 $X=1976698 $Y=881040
X87 6144 1 3 7643 7644 NOR2X4 $T=1981320 795760 1 180 $X=1976700 $Y=795358
X88 7666 1 3 7644 7494 NOR2X4 $T=1981320 815920 0 180 $X=1976700 $Y=810480
X89 7794 1 3 5901 7666 NOR2X4 $T=2003100 805840 1 0 $X=2003098 $Y=800400
X90 8521 1 3 8520 8162 NOR2X4 $T=2159520 876400 1 180 $X=2154900 $Y=875998
X91 2595 3 2592 2547 1 NAND2BX1 $T=939180 926800 0 180 $X=936540 $Y=921360
X92 3761 3 3743 3865 1 NAND2BX1 $T=1203840 785680 0 0 $X=1203838 $Y=785278
X93 5125 3 5029 5197 1 NAND2BX1 $T=1459920 836080 0 0 $X=1459918 $Y=835678
X94 5521 3 5523 5544 1 NAND2BX1 $T=1541100 856240 0 0 $X=1541098 $Y=855838
X95 5672 3 5539 5708 1 NAND2BX1 $T=1566180 785680 1 0 $X=1566178 $Y=780240
X96 168 3 169 5937 1 NAND2BX1 $T=1607760 745360 1 0 $X=1607758 $Y=739920
X97 343 3 218 217 1 NAND2BX1 $T=1789260 977200 1 180 $X=1786620 $Y=976798
X98 6942 3 6902 7013 1 NAND2BX1 $T=1839420 926800 0 0 $X=1839418 $Y=926398
X99 7227 3 7229 7214 1 NAND2BX1 $T=1892880 846160 1 180 $X=1890240 $Y=845758
X100 7301 3 7298 7315 1 NAND2BX1 $T=1910040 826000 1 0 $X=1910038 $Y=820560
X101 7493 3 7533 7481 1 NAND2BX1 $T=1955580 805840 0 180 $X=1952940 $Y=800400
X102 7666 3 7664 7652 1 NAND2BX1 $T=1983300 805840 1 180 $X=1980660 $Y=805438
X103 8179 3 8182 8121 1 NAND2BX1 $T=2091540 896560 1 180 $X=2088900 $Y=896158
X104 264 3 262 8390 1 NAND2BX1 $T=2141040 977200 1 180 $X=2138400 $Y=976798
X105 8682 3 8745 8681 1 NAND2BX1 $T=2211660 977200 0 180 $X=2209020 $Y=971760
X106 8897 3 8899 8835 1 NAND2BX1 $T=2240700 846160 0 180 $X=2238060 $Y=840720
X107 3391 3382 3 3362 1 3346 OAI21X1 $T=1116720 866320 1 180 $X=1113420 $Y=865918
X108 3476 3477 3 3456 1 3453 OAI21X1 $T=1137180 856240 1 180 $X=1133880 $Y=855838
X109 3800 3881 3 3791 1 3724 OAI21X1 $T=1200540 815920 1 180 $X=1197240 $Y=815518
X110 3741 3850 3 3791 1 3758 OAI21X1 $T=1204500 836080 1 0 $X=1204498 $Y=830640
X111 104 3967 3 4006 1 4110 OAI21X1 $T=1229580 957040 1 0 $X=1229578 $Y=951600
X112 4188 4213 3 4222 1 4232 OAI21X1 $T=1268520 755440 0 180 $X=1265220 $Y=750000
X113 5029 4957 3 5022 1 5028 OAI21X1 $T=1440120 826000 0 180 $X=1436820 $Y=820560
X114 4994 5154 3 5076 1 150 OAI21X1 $T=1461900 765520 1 180 $X=1458600 $Y=765118
X115 5516 5497 3 5474 1 5520 OAI21X1 $T=1537800 755440 0 0 $X=1537798 $Y=755038
X116 5937 5943 3 171 1 5938 OAI21X1 $T=1617000 745360 1 180 $X=1613700 $Y=744958
X117 226 7190 3 7215 1 7153 OAI21X1 $T=1888260 957040 0 0 $X=1888258 $Y=956638
X118 7388 7486 3 7426 1 7453 OAI21X1 $T=1947000 805840 1 180 $X=1943700 $Y=805438
X119 8384 8162 3 8413 1 8346 OAI21X1 $T=2135760 856240 0 0 $X=2135758 $Y=855838
X120 8616 8593 3 8629 1 8521 OAI21X1 $T=2180640 876400 0 0 $X=2180638 $Y=875998
X121 8836 8897 3 8899 1 8638 OAI21X1 $T=2238060 866320 1 0 $X=2238058 $Y=860880
X122 45 3 46 2397 1 47 OAI21XL $T=900240 967120 0 0 $X=900238 $Y=966718
X123 2546 3 46 2566 1 2567 OAI21XL $T=933240 946960 0 0 $X=933238 $Y=946558
X124 2594 3 46 2593 1 2548 OAI21XL $T=939840 926800 1 180 $X=937200 $Y=926398
X125 2595 3 2593 2592 1 2478 OAI21XL $T=947100 926800 1 180 $X=944460 $Y=926398
X126 2713 3 46 2735 1 2737 OAI21XL $T=961620 946960 0 0 $X=961618 $Y=946558
X127 2734 3 46 2736 1 2755 OAI21XL $T=962940 926800 0 0 $X=962938 $Y=926398
X128 2797 3 2800 2798 1 2778 OAI21XL $T=980100 926800 0 180 $X=977460 $Y=921360
X129 3320 3 3338 3340 1 3361 OAI21XL $T=1108140 846160 0 0 $X=1108138 $Y=845758
X130 3321 3 3345 3337 1 3339 OAI21XL $T=1112100 826000 0 180 $X=1109460 $Y=820560
X131 3343 3 80 3406 1 3507 OAI21XL $T=1125300 896560 1 0 $X=1125298 $Y=891120
X132 3461 3 3034 3475 1 3341 OAI21XL $T=1131900 836080 1 180 $X=1129260 $Y=835678
X133 3251 3 3455 3446 1 3448 OAI21XL $T=1135860 795760 0 180 $X=1133220 $Y=790320
X134 3478 3 3449 3460 1 3452 OAI21XL $T=1138500 916720 0 180 $X=1135860 $Y=911280
X135 3461 3 49 3475 1 3570 OAI21XL $T=1137180 836080 0 0 $X=1137178 $Y=835678
X136 84 3 71 3487 1 3520 OAI21XL $T=1145100 896560 0 0 $X=1145098 $Y=896158
X137 3478 3 86 3460 1 3593 OAI21XL $T=1147080 916720 0 0 $X=1147078 $Y=916318
X138 3479 3 3503 3506 1 3614 OAI21XL $T=1155000 775600 0 0 $X=1154998 $Y=775198
X139 3425 3 3034 3641 1 3506 OAI21XL $T=1160280 876400 1 180 $X=1157640 $Y=875998
X140 3457 3 3572 3592 1 3648 OAI21XL $T=1161600 846160 1 0 $X=1161598 $Y=840720
X141 76 3 86 49 1 3642 OAI21XL $T=1164240 926800 0 0 $X=1164238 $Y=926398
X142 3687 3 3670 3692 1 3711 OAI21XL $T=1176120 866320 0 0 $X=1176118 $Y=865918
X143 3668 3 3689 3693 1 3845 OAI21XL $T=1176120 946960 1 0 $X=1176118 $Y=941520
X144 3664 3 96 3704 1 3937 OAI21XL $T=1188000 977200 1 0 $X=1187998 $Y=971760
X145 3787 3 3573 3520 1 3785 OAI21XL $T=1198560 876400 0 180 $X=1195920 $Y=870960
X146 3665 3 100 3789 1 3787 OAI21XL $T=1199880 926800 0 180 $X=1197240 $Y=921360
X147 3845 3 3867 3593 1 3838 OAI21XL $T=1203840 916720 1 180 $X=1201200 $Y=916318
X148 3448 3 3848 3617 1 3797 OAI21XL $T=1206480 755440 1 180 $X=1203840 $Y=755038
X149 69 3 75 62 1 3878 OAI21XL $T=1206480 906640 0 0 $X=1206478 $Y=906238
X150 102 3 103 344 1 3885 OAI21XL $T=1210440 977200 0 0 $X=1210438 $Y=976798
X151 76 3 71 3878 1 3963 OAI21XL $T=1216380 906640 0 0 $X=1216378 $Y=906238
X152 3848 3 3849 3448 1 3951 OAI21XL $T=1223640 765520 1 180 $X=1221000 $Y=765118
X153 4077 3 4174 4186 1 4196 OAI21XL $T=1254660 775600 1 0 $X=1254658 $Y=770160
X154 4244 3 4233 4298 1 4414 OAI21XL $T=1281060 815920 0 0 $X=1281058 $Y=815518
X155 71 3 4307 65 1 4345 OAI21XL $T=1285020 866320 1 0 $X=1285018 $Y=860880
X156 5178 3 151 5173 1 5174 OAI21XL $T=1468500 745360 1 180 $X=1465860 $Y=744958
X157 5059 3 151 4994 1 5181 OAI21XL $T=1471800 775600 0 180 $X=1469160 $Y=770160
X158 5262 3 5278 5244 1 5264 OAI21XL $T=1492260 926800 0 180 $X=1489620 $Y=921360
X159 5315 3 5432 5278 1 5411 OAI21XL $T=1518000 926800 1 0 $X=1517998 $Y=921360
X160 5455 3 5733 5498 1 5754 OAI21XL $T=1574100 836080 1 0 $X=1574098 $Y=830640
X161 174 3 175 176 1 5981 OAI21XL $T=1618980 745360 1 0 $X=1618978 $Y=739920
X162 8161 3 8162 8178 1 8120 OAI21XL $T=2086260 876400 0 0 $X=2086258 $Y=875998
X163 8179 3 8178 8182 1 8139 OAI21XL $T=2094180 896560 0 0 $X=2094178 $Y=896158
X164 8283 3 8162 8269 1 8270 OAI21XL $T=2106720 866320 0 180 $X=2104080 $Y=860880
X165 8385 3 8324 8370 1 8267 OAI21XL $T=2132460 876400 0 180 $X=2129820 $Y=870960
X166 8589 3 260 8593 1 8573 OAI21XL $T=2172720 866320 1 0 $X=2172718 $Y=860880
X167 8746 3 8743 8741 1 8679 OAI21XL $T=2201760 886480 0 180 $X=2199120 $Y=881040
X168 271 3 8682 8745 1 8633 OAI21XL $T=2202420 977200 1 0 $X=2202418 $Y=971760
X169 5628 5767 5897 3 1 XOR2X4 $T=1574760 815920 0 0 $X=1574758 $Y=815518
X170 5896 5898 5932 3 1 XOR2X4 $T=1601820 946960 0 0 $X=1601818 $Y=946558
X171 5655 5914 6192 3 1 XOR2X4 $T=1610400 765520 1 0 $X=1610398 $Y=760080
X172 120 5961 6818 3 1 XOR2X4 $T=1768140 896560 0 0 $X=1768138 $Y=896158
X173 7424 7404 232 3 1 XOR2X4 $T=1938420 826000 1 180 $X=1927200 $Y=825598
X174 7481 7530 237 3 1 XOR2X4 $T=1946340 846160 0 0 $X=1946338 $Y=845758
X175 7552 7528 239 3 1 XOR2X4 $T=1958220 926800 1 0 $X=1958218 $Y=921360
X176 7652 7619 240 3 1 XOR2X4 $T=1983300 836080 1 180 $X=1972080 $Y=835678
X177 7616 7621 241 3 1 XOR2X4 $T=1973400 957040 0 0 $X=1973398 $Y=956638
X178 2367 3 1 2546 INVX1 $T=928620 946960 0 0 $X=928618 $Y=946558
X179 2478 3 1 2566 INVX1 $T=942480 946960 1 180 $X=941160 $Y=946558
X180 2735 3 1 2780 INVX1 $T=986040 946960 1 0 $X=986038 $Y=941520
X181 65 3 1 50 INVX1 $T=1039500 916720 0 180 $X=1038180 $Y=911280
X182 62 3 1 3155 INVX1 $T=1063260 896560 1 180 $X=1061940 $Y=896158
X183 3455 3 1 3475 INVX1 $T=1135200 815920 1 0 $X=1135198 $Y=810480
X184 3449 3 1 3487 INVX1 $T=1141140 896560 0 0 $X=1141138 $Y=896158
X185 3379 3 1 3503 INVX1 $T=1147080 785680 1 0 $X=1147078 $Y=780240
X186 3453 3 1 3572 INVX1 $T=1148400 846160 1 0 $X=1148398 $Y=840720
X187 3479 3 1 3623 INVX1 $T=1166220 785680 1 0 $X=1166218 $Y=780240
X188 3483 3 1 3689 INVX1 $T=1166220 946960 0 0 $X=1166218 $Y=946558
X189 3648 3 1 3720 INVX1 $T=1168860 846160 0 0 $X=1168858 $Y=845758
X190 3507 3 1 3670 INVX1 $T=1168860 886480 1 0 $X=1168858 $Y=881040
X191 3720 3 1 3725 INVX1 $T=1184040 846160 0 0 $X=1184038 $Y=845758
X192 3741 3 1 3842 INVX1 $T=1189980 826000 1 0 $X=1189978 $Y=820560
X193 3761 3 1 3764 INVX1 $T=1192620 785680 1 0 $X=1192618 $Y=780240
X194 3797 3 1 3802 INVX1 $T=1199880 765520 1 0 $X=1199878 $Y=760080
X195 3842 3 1 3800 INVX1 $T=1201860 805840 1 180 $X=1200540 $Y=805438
X196 3850 3 1 3882 INVX1 $T=1213740 836080 1 0 $X=1213738 $Y=830640
X197 3885 3 1 3967 INVX1 $T=1216380 957040 1 0 $X=1216378 $Y=951600
X198 3946 3 1 3875 INVX1 $T=1220340 836080 1 180 $X=1219020 $Y=835678
X199 4033 3 1 4049 INVX1 $T=1234200 896560 0 0 $X=1234198 $Y=896158
X200 3937 3 1 4091 INVX1 $T=1234200 967120 0 0 $X=1234198 $Y=966718
X201 4105 3 1 4130 INVX1 $T=1247400 936880 1 0 $X=1247398 $Y=931440
X202 4053 3 1 4169 INVX1 $T=1250040 886480 0 0 $X=1250038 $Y=886078
X203 4173 3 1 4312 INVX1 $T=1286340 926800 0 0 $X=1286338 $Y=926398
X204 4274 3 1 4476 INVX1 $T=1288980 977200 1 0 $X=1288978 $Y=971760
X205 4240 3 1 4324 INVX1 $T=1290960 795760 1 180 $X=1289640 $Y=795358
X206 4333 3 1 4417 INVX1 $T=1291620 896560 0 0 $X=1291618 $Y=896158
X207 4042 3 1 4416 INVX1 $T=1298880 775600 0 0 $X=1298878 $Y=775198
X208 4085 3 1 4439 INVX1 $T=1302180 846160 0 0 $X=1302178 $Y=845758
X209 4436 3 1 4415 INVX1 $T=1303500 745360 0 180 $X=1302180 $Y=739920
X210 3952 3 1 4715 INVX1 $T=1312740 815920 0 0 $X=1312738 $Y=815518
X211 4122 3 1 4581 INVX1 $T=1320660 795760 1 0 $X=1320658 $Y=790320
X212 3980 3 1 4582 INVX1 $T=1320660 876400 1 0 $X=1320658 $Y=870960
X213 5006 3 1 5050 INVX1 $T=1432860 775600 1 0 $X=1432858 $Y=770160
X214 4993 3 1 149 INVX1 $T=1448700 745360 0 0 $X=1448698 $Y=744958
X215 5039 3 1 5117 INVX1 $T=1448700 785680 1 0 $X=1448698 $Y=780240
X216 5053 3 1 5134 INVX1 $T=1453980 785680 0 0 $X=1453978 $Y=785278
X217 5125 3 1 5137 INVX1 $T=1456620 826000 0 0 $X=1456618 $Y=825598
X218 5059 3 1 5136 INVX1 $T=1464540 775600 0 0 $X=1464538 $Y=775198
X219 5198 3 1 5238 INVX1 $T=1475100 866320 0 0 $X=1475098 $Y=865918
X220 5176 3 1 5243 INVX1 $T=1477740 876400 1 0 $X=1477738 $Y=870960
X221 150 3 1 5314 INVX1 $T=1481040 765520 0 0 $X=1481038 $Y=765118
X222 152 3 1 5311 INVX1 $T=1496220 795760 1 0 $X=1496218 $Y=790320
X223 5319 3 1 5432 INVX1 $T=1511400 926800 1 0 $X=1511398 $Y=921360
X224 5298 3 1 161 INVX1 $T=1524600 967120 0 0 $X=1524598 $Y=966718
X225 5625 3 1 5675 INVX1 $T=1556280 886480 0 0 $X=1556278 $Y=886078
X226 5589 3 1 5733 INVX1 $T=1570140 836080 1 0 $X=1570138 $Y=830640
X227 5413 3 1 5758 INVX1 $T=1574760 755440 1 0 $X=1574758 $Y=750000
X228 5455 3 1 5774 INVX1 $T=1576740 846160 1 0 $X=1576738 $Y=840720
X229 5581 3 1 5760 INVX1 $T=1579380 916720 0 0 $X=1579378 $Y=916318
X230 5656 3 1 5761 INVX1 $T=1585980 957040 0 180 $X=1584660 $Y=951600
X231 5787 3 1 5833 INVX1 $T=1587300 775600 0 0 $X=1587298 $Y=775198
X232 6059 3 1 6035 INVX1 $T=1644060 936880 1 0 $X=1644058 $Y=931440
X233 5936 3 1 192 INVX1 $T=1644720 755440 0 0 $X=1644718 $Y=755038
X234 6067 3 1 6077 INVX1 $T=1645380 946960 1 0 $X=1645378 $Y=941520
X235 6126 3 1 6091 INVX1 $T=1656600 916720 1 180 $X=1655280 $Y=916318
X236 6207 3 1 6161 INVX1 $T=1676400 967120 1 0 $X=1676398 $Y=961680
X237 6226 3 1 6194 INVX1 $T=1679040 926800 1 0 $X=1679038 $Y=921360
X238 6420 3 1 6423 INVX1 $T=1716660 957040 0 0 $X=1716658 $Y=956638
X239 6422 3 1 6426 INVX1 $T=1717980 926800 1 0 $X=1717978 $Y=921360
X240 6405 3 1 6462 INVX1 $T=1728540 946960 0 0 $X=1728538 $Y=946558
X241 7061 3 1 7081 INVX1 $T=1849320 957040 0 0 $X=1849318 $Y=956638
X242 7084 3 1 7106 INVX1 $T=1860540 886480 0 0 $X=1860538 $Y=886078
X243 7080 3 1 6991 INVX1 $T=1863840 936880 0 180 $X=1862520 $Y=931440
X244 7190 3 1 7177 INVX1 $T=1882980 957040 0 0 $X=1882978 $Y=956638
X245 7192 3 1 7154 INVX1 $T=1884300 866320 1 180 $X=1882980 $Y=865918
X246 7213 3 1 7235 INVX1 $T=1888260 896560 1 0 $X=1888258 $Y=891120
X247 7388 3 1 7386 INVX1 $T=1928520 805840 1 180 $X=1927200 $Y=805438
X248 7408 3 1 7412 INVX1 $T=1932480 886480 0 0 $X=1932478 $Y=886078
X249 7482 3 1 7490 INVX1 $T=1948320 916720 0 0 $X=1948318 $Y=916318
X250 7644 3 1 7697 INVX1 $T=1987920 815920 0 0 $X=1987918 $Y=815518
X251 7717 3 1 7684 INVX1 $T=1998480 826000 0 0 $X=1998478 $Y=825598
X252 7907 3 1 7838 INVX1 $T=2032140 906640 0 0 $X=2032138 $Y=906238
X253 7939 3 1 7897 INVX1 $T=2036100 836080 1 180 $X=2034780 $Y=835678
X254 7996 3 1 7853 INVX1 $T=2046660 876400 0 180 $X=2045340 $Y=870960
X255 7997 3 1 7979 INVX1 $T=2049960 957040 1 0 $X=2049958 $Y=951600
X256 8112 3 1 7926 INVX1 $T=2067120 826000 0 180 $X=2065800 $Y=820560
X257 8003 3 1 8073 INVX1 $T=2069760 846160 0 180 $X=2068440 $Y=840720
X258 8095 3 1 8110 INVX1 $T=2071080 896560 0 0 $X=2071078 $Y=896158
X259 7941 3 1 8138 INVX1 $T=2073720 805840 0 0 $X=2073718 $Y=805438
X260 8162 3 1 8140 INVX1 $T=2082960 886480 1 180 $X=2081640 $Y=886078
X261 8141 3 1 8146 INVX1 $T=2092200 815920 1 0 $X=2092198 $Y=810480
X262 8266 3 1 8111 INVX1 $T=2096160 826000 0 180 $X=2094840 $Y=820560
X263 8305 3 1 8283 INVX1 $T=2109360 866320 0 180 $X=2108040 $Y=860880
X264 8325 3 1 8327 INVX1 $T=2117280 846160 1 180 $X=2115960 $Y=845758
X265 259 3 1 263 INVX1 $T=2137740 967120 1 0 $X=2137738 $Y=961680
X266 8458 3 1 8388 INVX1 $T=2143020 876400 1 180 $X=2141700 $Y=875998
X267 8385 3 1 8417 INVX1 $T=2145660 866320 0 180 $X=2144340 $Y=860880
X268 8499 3 1 8500 INVX1 $T=2150940 977200 0 180 $X=2149620 $Y=971760
X269 268 3 1 8502 INVX1 $T=2156220 977200 0 180 $X=2154900 $Y=971760
X270 8572 3 1 8547 INVX1 $T=2170080 876400 1 180 $X=2168760 $Y=875998
X271 8589 3 1 8632 INVX1 $T=2181300 866320 1 0 $X=2181298 $Y=860880
X272 272 3 1 255 INVX1 $T=2184600 946960 0 180 $X=2183280 $Y=941520
X273 8761 3 1 8659 INVX1 $T=2195820 856240 1 180 $X=2194500 $Y=855838
X274 8758 3 1 8850 INVX1 $T=2233440 866320 0 0 $X=2233438 $Y=865918
X275 63 78 1 3319 3382 3 AOI21X2 $T=1120680 957040 0 180 $X=1116060 $Y=951600
X276 155 5219 1 5160 5214 3 AOI21X2 $T=1480380 846160 1 180 $X=1475760 $Y=845758
X277 155 5238 1 5243 5293 3 AOI21X2 $T=1483680 876400 1 0 $X=1483678 $Y=870960
X278 5260 155 1 5297 5362 3 AOI21X2 $T=1492920 745360 0 0 $X=1492918 $Y=744958
X279 5326 5319 1 5264 5301 3 AOI21X2 $T=1500180 926800 0 180 $X=1495560 $Y=921360
X280 160 5379 1 5319 5406 3 AOI21X2 $T=1513380 957040 0 180 $X=1508760 $Y=951600
X281 5688 5675 1 5629 5685 3 AOI21X2 $T=1568160 886480 1 180 $X=1563540 $Y=886078
X282 5712 5716 1 5520 5727 3 AOI21X2 $T=1573440 765520 0 180 $X=1568820 $Y=760080
X283 5768 5717 1 5761 5756 3 AOI21X2 $T=1582680 967120 0 180 $X=1578060 $Y=961680
X284 5688 5709 1 5754 5767 3 AOI21X2 $T=1579380 836080 1 0 $X=1579378 $Y=830640
X285 6069 181 1 5981 6068 3 AOI21X2 $T=1646700 745360 1 180 $X=1642080 $Y=744958
X286 7108 7153 1 7081 7147 3 AOI21X2 $T=1874400 957040 1 180 $X=1869780 $Y=956638
X287 7489 7527 1 7453 7530 3 AOI21X2 $T=1952940 836080 1 180 $X=1948320 $Y=835678
X288 7527 7697 1 7684 7619 3 AOI21X2 $T=1989900 826000 1 180 $X=1985280 $Y=825598
X289 1 2595 2594 2367 3 NOR2X1 $T=939180 936880 1 180 $X=937200 $Y=936478
X290 1 2695 2615 2595 3 NOR2X1 $T=952380 916720 1 180 $X=950400 $Y=916318
X291 1 2797 2820 2779 3 NOR2X1 $T=982080 926800 1 180 $X=980100 $Y=926398
X292 1 2841 2825 2797 3 NOR2X1 $T=986040 906640 1 180 $X=984060 $Y=906238
X293 1 2865 2864 2820 3 NOR2X1 $T=1005840 926800 1 180 $X=1003860 $Y=926398
X294 1 63 78 3319 3 NOR2X1 $T=1111440 957040 1 0 $X=1111438 $Y=951600
X295 1 79 62 3449 3 NOR2X1 $T=1126620 977200 1 0 $X=1126618 $Y=971760
X296 1 74 65 3455 3 NOR2X1 $T=1136520 826000 1 180 $X=1134540 $Y=825598
X297 1 84 3449 3425 3 NOR2X1 $T=1138500 896560 1 180 $X=1136520 $Y=896158
X298 1 3035 72 3478 3 NOR2X1 $T=1149720 906640 0 180 $X=1147740 $Y=901200
X299 1 3424 3361 3741 3 NOR2X1 $T=1167540 826000 0 0 $X=1167538 $Y=825598
X300 1 3717 3711 3761 3 NOR2X1 $T=1189320 785680 0 0 $X=1189318 $Y=785278
X301 1 3915 3908 4053 3 NOR2X1 $T=1215720 896560 1 0 $X=1215718 $Y=891120
X302 1 3844 3801 3946 3 NOR2X1 $T=1218360 846160 1 0 $X=1218358 $Y=840720
X303 1 4047 4091 4033 3 NOR2X1 $T=1244760 916720 0 0 $X=1244758 $Y=916318
X304 1 109 4080 4132 3 NOR2X1 $T=1247400 967120 1 0 $X=1247398 $Y=961680
X305 1 4194 4196 4213 3 NOR2X1 $T=1258620 755440 0 0 $X=1258618 $Y=755038
X306 1 4359 4414 4438 3 NOR2X1 $T=1307460 755440 0 0 $X=1307458 $Y=755038
X307 1 4944 4947 4957 3 NOR2X1 $T=1421640 826000 0 180 $X=1419660 $Y=820560
X308 1 4981 4921 5059 3 NOR2X1 $T=1425600 785680 1 0 $X=1425598 $Y=780240
X309 1 5175 5123 5198 3 NOR2X1 $T=1466520 866320 0 0 $X=1466518 $Y=865918
X310 1 5059 5154 153 3 NOR2X1 $T=1471140 765520 0 0 $X=1471138 $Y=765118
X311 1 5059 152 5221 3 NOR2X1 $T=1472460 785680 1 0 $X=1472458 $Y=780240
X312 1 5078 5198 5219 3 NOR2X1 $T=1472460 856240 1 0 $X=1472458 $Y=850800
X313 1 5178 152 5213 3 NOR2X1 $T=1474440 755440 1 0 $X=1474438 $Y=750000
X314 1 156 5203 5298 3 NOR2X1 $T=1488300 977200 0 0 $X=1488298 $Y=976798
X315 1 5581 5679 5728 3 NOR2X1 $T=1569480 916720 1 0 $X=1569478 $Y=911280
X316 1 5937 5936 5934 3 NOR2X1 $T=1615020 775600 0 180 $X=1613040 $Y=770160
X317 1 5932 7234 7190 3 NOR2X1 $T=1892880 957040 1 0 $X=1892878 $Y=951600
X318 1 8179 8161 8142 3 NOR2X1 $T=2083620 896560 1 180 $X=2081640 $Y=896158
X319 1 8445 8462 8325 3 NOR2X1 $T=2148960 866320 1 180 $X=2146980 $Y=865918
X320 1 8616 8589 8572 3 NOR2X1 $T=2174700 876400 1 180 $X=2172720 $Y=875998
X321 1 273 8682 8612 3 NOR2X1 $T=2195820 967120 0 0 $X=2195818 $Y=966718
X322 1 8791 8698 8743 3 NOR2X1 $T=2203740 896560 1 180 $X=2201760 $Y=896158
X323 1 8758 8743 8674 3 NOR2X1 $T=2206380 876400 1 180 $X=2204400 $Y=875998
X324 1 8859 8914 8897 3 NOR2X1 $T=2245320 876400 1 0 $X=2245318 $Y=870960
X325 1 8860 8943 8878 3 NOR2X1 $T=2254560 876400 0 180 $X=2252580 $Y=870960
X326 3455 3461 3 1 3379 NOR2X2 $T=1140480 826000 1 180 $X=1137180 $Y=825598
X327 4968 5023 3 1 5125 NOR2X2 $T=1444080 836080 0 0 $X=1444078 $Y=835678
X328 5116 5055 3 1 5078 NOR2X2 $T=1451340 856240 1 180 $X=1448040 $Y=855838
X329 5125 4957 3 1 5135 NOR2X2 $T=1453320 826000 1 0 $X=1453318 $Y=820560
X330 5118 5008 3 1 5294 NOR2X2 $T=1479720 967120 1 0 $X=1479718 $Y=961680
X331 5220 5163 3 1 5262 NOR2X2 $T=1482360 926800 1 0 $X=1482358 $Y=921360
X332 5282 5072 3 1 5315 NOR2X2 $T=1490940 936880 0 0 $X=1490938 $Y=936478
X333 5262 5315 3 1 5326 NOR2X2 $T=1503480 926800 1 0 $X=1503478 $Y=921360
X334 5298 5294 3 1 5379 NOR2X2 $T=1503480 967120 1 0 $X=1503478 $Y=961680
X335 5429 4193 3 1 5413 NOR2X2 $T=1519980 755440 0 180 $X=1516680 $Y=750000
X336 5430 4439 3 1 5521 NOR2X2 $T=1519980 856240 1 180 $X=1516680 $Y=855838
X337 5364 4715 3 1 5455 NOR2X2 $T=1522620 826000 0 0 $X=1522618 $Y=825598
X338 5400 4452 3 1 5513 NOR2X2 $T=1523940 815920 0 0 $X=1523938 $Y=815518
X339 5401 4582 3 1 5625 NOR2X2 $T=1529220 876400 1 0 $X=1529218 $Y=870960
X340 162 4494 3 1 5497 NOR2X2 $T=1532520 745360 0 0 $X=1532518 $Y=744958
X341 5547 4312 3 1 5581 NOR2X2 $T=1545720 926800 1 0 $X=1545718 $Y=921360
X342 5402 4417 3 1 5679 NOR2X2 $T=1553640 906640 1 180 $X=1550340 $Y=906238
X343 5267 4581 3 1 5649 NOR2X2 $T=1561560 795760 0 180 $X=1558260 $Y=790320
X344 5413 5497 3 1 5712 NOR2X2 $T=1560900 755440 0 0 $X=1560898 $Y=755038
X345 5672 5649 3 1 5787 NOR2X2 $T=1578720 785680 1 0 $X=1578718 $Y=780240
X346 178 208 3 1 6050 NOR2X2 $T=1698180 896560 0 180 $X=1694880 $Y=891120
X347 209 178 3 1 6066 NOR2X2 $T=1697520 916720 1 0 $X=1697518 $Y=911280
X348 5963 6901 3 1 6898 NOR2X2 $T=1823580 906640 1 180 $X=1820280 $Y=906238
X349 6927 5939 3 1 6942 NOR2X2 $T=1833480 936880 0 180 $X=1830180 $Y=931440
X350 6898 6942 3 1 7062 NOR2X2 $T=1838760 916720 1 0 $X=1838758 $Y=911280
X351 7232 5897 3 1 7227 NOR2X2 $T=1893540 826000 0 180 $X=1890240 $Y=820560
X352 7301 7227 3 1 7300 NOR2X2 $T=1900800 826000 0 0 $X=1900798 $Y=825598
X353 7317 6193 3 1 7301 NOR2X2 $T=1904100 815920 0 180 $X=1900800 $Y=810480
X354 7405 231 3 1 7375 NOR2X2 $T=1927860 876400 0 180 $X=1924560 $Y=870960
X355 6192 7410 3 1 7388 NOR2X2 $T=1929180 785680 1 180 $X=1925880 $Y=785278
X356 7446 233 3 1 7428 NOR2X2 $T=1939740 866320 1 0 $X=1939738 $Y=860880
X357 7598 7484 3 1 7611 NOR2X2 $T=1969440 886480 1 0 $X=1969438 $Y=881040
X358 7640 6818 3 1 7622 NOR2X2 $T=1976700 926800 0 0 $X=1976698 $Y=926398
X359 8092 8141 3 1 8050 NOR2X2 $T=2080980 826000 1 0 $X=2080978 $Y=820560
X360 266 264 3 1 8499 NOR2X2 $T=2148960 977200 0 0 $X=2148958 $Y=976798
X361 8547 260 3 1 8520 NOR2X2 $T=2162820 876400 0 0 $X=2162818 $Y=875998
X362 8810 278 3 1 8682 NOR2X2 $T=2215620 977200 0 0 $X=2215618 $Y=976798
X363 8792 8851 3 1 8758 NOR2X2 $T=2228160 876400 1 180 $X=2224860 $Y=875998
X364 8878 8897 3 1 8657 NOR2X2 $T=2233440 876400 0 180 $X=2230140 $Y=870960
X365 3155 4240 3 1 4418 OR2XL $T=1298880 785680 1 0 $X=1298878 $Y=780240
X366 8282 258 3 1 8117 OR2XL $T=2106060 906640 1 180 $X=2103420 $Y=906238
X367 3720 3381 3763 3 1 NAND2X2 $T=1195920 846160 1 180 $X=1192620 $Y=845758
X368 5219 5135 152 3 1 NAND2X2 $T=1476420 815920 0 0 $X=1476418 $Y=815518
X369 4476 163 164 3 1 NAND2X2 $T=1540440 977200 1 180 $X=1537140 $Y=976798
X370 5401 4582 5538 3 1 NAND2X2 $T=1545060 876400 0 180 $X=1541760 $Y=870960
X371 5410 4416 5539 3 1 NAND2X2 $T=1546380 775600 1 180 $X=1543080 $Y=775198
X372 5712 5787 5936 3 1 NAND2X2 $T=1595220 775600 0 180 $X=1591920 $Y=770160
X373 195 191 6125 3 1 NAND2X2 $T=1653300 745360 1 0 $X=1653298 $Y=739920
X374 6927 5939 6902 3 1 NAND2X2 $T=1825560 936880 0 180 $X=1822260 $Y=931440
X375 7083 7085 7082 3 1 NAND2X2 $T=1859220 876400 0 180 $X=1855920 $Y=870960
X376 5966 7150 7151 3 1 NAND2X2 $T=1871760 876400 0 0 $X=1871758 $Y=875998
X377 7232 5897 7229 3 1 NAND2X2 $T=1894200 815920 1 180 $X=1890900 $Y=815518
X378 7237 7257 229 3 1 NAND2X2 $T=1898160 906640 0 0 $X=1898158 $Y=906238
X379 5965 7238 226 3 1 NAND2X2 $T=1904760 977200 0 180 $X=1901460 $Y=971760
X380 7386 7426 7424 3 1 NAND2X2 $T=1935120 805840 1 180 $X=1931820 $Y=805438
X381 7405 231 7408 3 1 NAND2X2 $T=1932480 876400 1 0 $X=1932478 $Y=870960
X382 6192 7410 7426 3 1 NAND2X2 $T=1935780 795760 1 0 $X=1935778 $Y=790320
X383 7427 7482 7484 3 1 NAND2X2 $T=1949640 886480 0 180 $X=1946340 $Y=881040
X384 7482 7454 7552 3 1 NAND2X2 $T=1947660 906640 0 0 $X=1947658 $Y=906238
X385 7526 7494 7551 3 1 NAND2X2 $T=1959540 815920 1 180 $X=1956240 $Y=815518
X386 7637 6273 7620 3 1 NAND2X2 $T=1976040 876400 0 0 $X=1976038 $Y=875998
X387 7640 6818 7649 3 1 NAND2X2 $T=1977360 926800 1 0 $X=1977358 $Y=921360
X388 7794 5901 7664 3 1 NAND2X2 $T=1999800 805840 0 0 $X=1999798 $Y=805438
X389 7810 7834 7997 3 1 NAND2X2 $T=2029500 957040 0 0 $X=2029498 $Y=956638
X390 247 7877 7908 3 1 NAND2X2 $T=2033460 936880 1 180 $X=2030160 $Y=936478
X391 8499 8612 8589 3 1 NAND2X2 $T=2176020 967120 1 180 $X=2172720 $Y=966718
X392 5160 1 5135 5028 3 151 AOI21X4 $T=1465860 815920 1 180 $X=1459260 $Y=815518
X393 5540 1 5589 5586 3 5580 AOI21X4 $T=1554960 836080 0 180 $X=1548360 $Y=830640
X394 5688 1 5590 5589 3 5755 AOI21X4 $T=1564200 856240 1 0 $X=1564198 $Y=850800
X395 5731 1 5728 5682 3 5678 AOI21X4 $T=1575420 926800 0 180 $X=1568820 $Y=921360
X396 5815 1 5548 5768 3 5898 AOI21X4 $T=1589940 967120 0 0 $X=1589938 $Y=966718
X397 5934 1 5677 5938 3 5961 AOI21X4 $T=1611060 785680 0 0 $X=1611058 $Y=785278
X398 7080 1 7062 6944 3 7084 AOI21X4 $T=1853280 916720 1 0 $X=1853278 $Y=911280
X399 7175 1 7083 7154 3 7105 AOI21X4 $T=1879020 866320 1 180 $X=1872420 $Y=865918
X400 7149 1 7300 7302 3 7303 AOI21X4 $T=1898820 836080 0 0 $X=1898818 $Y=835678
X401 7427 1 7429 7412 3 7422 AOI21X4 $T=1942380 886480 1 180 $X=1935780 $Y=886078
X402 7527 1 7494 7480 3 7404 AOI21X4 $T=1952280 826000 0 180 $X=1945680 $Y=820560
X403 7526 1 7480 7570 3 7573 AOI21X4 $T=1956900 815920 1 0 $X=1956898 $Y=810480
X404 7611 1 7577 7618 3 7621 AOI21X4 $T=1970100 896560 0 0 $X=1970098 $Y=896158
X405 8612 1 268 8633 3 8593 AOI21X4 $T=2179320 967120 0 0 $X=2179318 $Y=966718
X406 3706 1 3727 3 3747 AND2X2 $T=1184700 826000 1 0 $X=1184698 $Y=820560
X407 4062 1 4050 3 4071 AND2X2 $T=1238820 856240 1 0 $X=1238818 $Y=850800
X408 4169 1 4139 3 4063 AND2X2 $T=1249380 866320 1 180 $X=1246740 $Y=865918
X409 4032 1 4169 3 4187 AND2X2 $T=1255980 886480 0 0 $X=1255978 $Y=886078
X410 5136 1 4994 3 5179 AND2X2 $T=1466520 795760 1 0 $X=1466518 $Y=790320
X411 5577 1 5474 3 5655 AND2X2 $T=1548360 755440 0 0 $X=1548358 $Y=755038
X412 5548 1 164 3 345 AND2X2 $T=1591920 977200 0 0 $X=1591918 $Y=976798
X413 7941 1 7971 3 8089 AND2X2 $T=2065140 815920 1 0 $X=2065138 $Y=810480
X414 5301 3 5358 1 155 NAND2X4 $T=1498200 906640 0 0 $X=1498198 $Y=906238
X415 5540 3 5590 1 5673 NAND2X4 $T=1558260 836080 1 0 $X=1558258 $Y=830640
X416 4581 3 5267 1 5729 NAND2X4 $T=1566180 795760 1 0 $X=1566178 $Y=790320
X417 233 3 7446 1 7454 NAND2X4 $T=1940400 866320 0 0 $X=1940398 $Y=865918
X418 6144 3 7643 1 7717 NAND2X4 $T=1991220 795760 0 0 $X=1991218 $Y=795358
X419 7881 3 7895 1 7148 NAND2X4 $T=2024220 856240 1 0 $X=2024218 $Y=850800
X420 8266 3 7975 1 8004 NAND2X4 $T=2101440 815920 0 0 $X=2101438 $Y=815518
X421 2505 2504 3 1 2366 OR2X2 $T=922680 946960 1 180 $X=920040 $Y=946558
X422 2886 2884 3 1 2712 OR2X2 $T=998580 946960 0 180 $X=995940 $Y=941520
X423 63 49 3 1 3460 OR2X2 $T=1145760 916720 0 180 $X=1143120 $Y=911280
X424 3758 3661 3 1 3691 OR2X2 $T=1182720 836080 0 180 $X=1180080 $Y=830640
X425 3339 3661 3 1 3719 OR2X2 $T=1181400 826000 1 0 $X=1181398 $Y=820560
X426 3936 4110 3 1 4113 OR2X2 $T=1255980 946960 0 0 $X=1255978 $Y=946558
X427 4276 4273 3 1 4262 OR2X2 $T=1278420 775600 1 180 $X=1275780 $Y=775198
X428 115 116 3 1 4561 OR2X2 $T=1337160 936880 1 0 $X=1337158 $Y=931440
X429 4987 4984 3 1 148 OR2X2 $T=1430220 745360 0 0 $X=1430218 $Y=744958
X430 4923 4966 3 1 5053 OR2X2 $T=1432860 785680 0 0 $X=1432858 $Y=785278
X431 4958 5038 3 1 5069 OR2X2 $T=1442760 775600 1 0 $X=1442758 $Y=770160
X432 5320 158 3 1 5358 OR2X2 $T=1498860 946960 1 0 $X=1498858 $Y=941520
X433 5627 4453 3 1 5717 OR2X2 $T=1561560 957040 1 0 $X=1561558 $Y=951600
X434 7102 5964 3 1 7108 OR2X2 $T=1861860 957040 1 0 $X=1861858 $Y=951600
X435 5965 7238 3 1 224 OR2X2 $T=1896180 977200 0 180 $X=1893540 $Y=971760
X436 7667 6668 3 1 7723 OR2X2 $T=1992540 916720 0 0 $X=1992538 $Y=916318
X437 7838 7836 3 1 7667 OR2X2 $T=2014320 916720 1 180 $X=2011680 $Y=916318
X438 245 246 3 1 7810 OR2X2 $T=2013660 977200 0 0 $X=2013658 $Y=976798
X439 7924 7896 3 1 7907 OR2X2 $T=2032800 896560 0 180 $X=2030160 $Y=891120
X440 8004 8072 3 1 8057 OR2X2 $T=2073060 836080 1 180 $X=2070420 $Y=835678
X441 8264 8207 3 1 8268 OR2X2 $T=2102100 886480 1 0 $X=2102098 $Y=881040
X442 8326 8328 3 1 8387 OR2X2 $T=2117940 896560 1 0 $X=2117938 $Y=891120
X443 8443 8389 3 1 8393 OR2X2 $T=2143680 886480 1 180 $X=2141040 $Y=886078
X444 2366 3 1 2367 45 NAND2XL $T=894300 946960 0 0 $X=894298 $Y=946558
X445 2712 3 1 2779 2594 NAND2XL $T=958980 936880 0 180 $X=957000 $Y=931440
X446 2735 3 1 2712 2640 NAND2XL $T=970860 946960 1 180 $X=968880 $Y=946558
X447 2865 3 1 2864 2800 NAND2XL $T=1012440 926800 1 180 $X=1010460 $Y=926398
X448 3758 3 1 3661 3727 NAND2XL $T=1193940 836080 0 180 $X=1191960 $Y=830640
X449 3791 3 1 3842 3918 NAND2XL $T=1207140 815920 1 0 $X=1207138 $Y=810480
X450 3908 3 1 3915 4032 NAND2XL $T=1213080 886480 0 0 $X=1213078 $Y=886078
X451 3801 3 1 3844 4050 NAND2XL $T=1218360 856240 1 0 $X=1218358 $Y=850800
X452 3875 3 1 3872 4062 NAND2XL $T=1226280 836080 0 0 $X=1226278 $Y=835678
X453 4196 3 1 4194 4222 NAND2XL $T=1268520 755440 1 180 $X=1266540 $Y=755038
X454 3155 3 1 4240 4273 NAND2XL $T=1280400 785680 1 180 $X=1278420 $Y=785278
X455 89 3 1 49 4240 NAND2XL $T=1282380 836080 1 0 $X=1282378 $Y=830640
X456 5038 3 1 4958 5006 NAND2XL $T=1440780 775600 0 0 $X=1440778 $Y=775198
X457 4993 3 1 148 5071 NAND2XL $T=1442100 745360 0 0 $X=1442098 $Y=744958
X458 5516 3 1 5758 5831 NAND2XL $T=1582020 765520 0 0 $X=1582018 $Y=765118
X459 7108 3 1 7061 7103 NAND2XL $T=1866480 957040 1 180 $X=1864500 $Y=956638
X460 7151 3 1 7085 7152 NAND2XL $T=1877700 876400 0 0 $X=1877698 $Y=875998
X461 7192 3 1 7083 7233 NAND2XL $T=1888260 876400 1 0 $X=1888258 $Y=870960
X462 8218 3 1 255 8182 NAND2XL $T=2102100 926800 1 180 $X=2100120 $Y=926398
X463 258 3 1 8282 8122 NAND2XL $T=2105400 916720 0 180 $X=2103420 $Y=911280
X464 8328 3 1 8326 8350 NAND2XL $T=2120580 886480 0 0 $X=2120578 $Y=886078
X465 8350 3 1 8387 8347 NAND2XL $T=2122560 876400 1 180 $X=2120580 $Y=875998
X466 8393 3 1 8327 8384 NAND2XL $T=2127840 856240 1 180 $X=2125860 $Y=855838
X467 8458 3 1 8393 8412 NAND2XL $T=2148960 856240 1 180 $X=2146980 $Y=855838
X468 8791 3 1 8698 8741 NAND2XL $T=2220240 896560 0 0 $X=2220238 $Y=896158
X469 8829 3 1 8632 8812 NAND2XL $T=2222220 856240 1 180 $X=2220240 $Y=855838
X470 65 89 3 1 INVX4 $T=1154340 815920 0 0 $X=1154338 $Y=815518
X471 5678 5688 3 1 INVX4 $T=1568820 866320 1 0 $X=1568818 $Y=860880
X472 5727 181 3 1 INVX4 $T=1628880 755440 0 0 $X=1628878 $Y=755038
X473 222 223 3 1 INVX4 $T=1874400 977200 0 180 $X=1871760 $Y=971760
X474 7977 7904 3 1 INVX4 $T=2067780 926800 0 0 $X=2067778 $Y=926398
X475 2780 2779 1 2778 2593 3 AOI21X1 $T=974820 926800 1 180 $X=972180 $Y=926398
X476 3428 3388 1 3389 3345 3 AOI21X1 $T=1122660 936880 1 180 $X=1120020 $Y=936478
X477 3617 3847 1 3849 3871 3 AOI21X1 $T=1203840 765520 0 0 $X=1203838 $Y=765118
X478 108 4172 1 4132 4219 3 AOI21X1 $T=1267860 957040 0 180 $X=1265220 $Y=951600
X479 5117 5069 1 5050 5076 3 AOI21X1 $T=1450680 775600 0 180 $X=1448040 $Y=770160
X480 148 150 1 149 5173 3 AOI21X1 $T=1461240 745360 0 0 $X=1461238 $Y=744958
X481 155 5213 1 5174 154 3 AOI21X1 $T=1477080 745360 0 180 $X=1474440 $Y=739920
X482 155 5200 1 5159 5215 3 AOI21X1 $T=1477740 785680 1 180 $X=1475100 $Y=785278
X483 155 5221 1 5181 5218 3 AOI21X1 $T=1479720 775600 1 180 $X=1477080 $Y=775198
X484 5239 155 1 5222 5248 3 AOI21X1 $T=1486320 826000 1 0 $X=1486318 $Y=820560
X485 5311 155 1 5318 5360 3 AOI21X1 $T=1501500 795760 1 0 $X=1501498 $Y=790320
X486 5407 160 1 5411 5405 3 AOI21X1 $T=1514700 936880 0 0 $X=1514698 $Y=936478
X487 5716 5758 1 5773 5895 3 AOI21X1 $T=1589280 755440 0 0 $X=1589278 $Y=755038
X488 7085 7106 1 7175 7213 3 AOI21X1 $T=1877040 886480 0 0 $X=1877038 $Y=886078
X489 8140 8142 1 8139 8095 3 AOI21X1 $T=2080980 896560 1 180 $X=2078340 $Y=896158
X490 8393 8417 1 8388 8413 3 AOI21X1 $T=2139720 866320 0 180 $X=2137080 $Y=860880
X491 8657 8640 1 8638 8634 3 AOI21X1 $T=2188560 866320 0 180 $X=2185920 $Y=860880
X492 8674 8638 1 8679 8629 3 AOI21X1 $T=2193840 876400 0 0 $X=2193838 $Y=875998
X493 8766 8640 1 8786 8782 3 AOI21X1 $T=2209680 866320 1 0 $X=2209678 $Y=860880
X494 8829 8640 1 8856 8828 3 AOI21X1 $T=2227500 856240 0 0 $X=2227498 $Y=855838
X495 4381 4438 3 4436 1 114 OAI21X2 $T=1313400 745360 0 180 $X=1308120 $Y=739920
X496 5176 5078 3 5161 1 5160 OAI21X2 $T=1469160 856240 0 180 $X=1463880 $Y=850800
X497 157 5294 3 5302 1 5319 OAI21X2 $T=1500840 967120 0 180 $X=1495560 $Y=961680
X498 5513 5498 3 5452 1 5586 OAI21X2 $T=1542420 826000 1 180 $X=1537140 $Y=825598
X499 5680 5679 3 5674 1 5682 OAI21X2 $T=1566180 916720 1 180 $X=1560900 $Y=916318
X500 6902 6898 3 6900 1 6944 OAI21X2 $T=1834140 916720 0 180 $X=1828860 $Y=911280
X501 6942 6991 3 6902 1 6948 OAI21X2 $T=1842720 936880 0 180 $X=1837440 $Y=931440
X502 7229 7301 3 7298 1 7302 OAI21X2 $T=1904100 815920 1 180 $X=1898820 $Y=815518
X503 7227 7258 3 7229 1 7335 OAI21X2 $T=1900800 846160 0 0 $X=1900798 $Y=845758
X504 7426 7493 3 7533 1 7570 OAI21X2 $T=1958220 805840 1 0 $X=1958218 $Y=800400
X505 7528 7484 3 7422 1 7574 OAI21X2 $T=1964820 896560 0 180 $X=1959540 $Y=891120
X506 7422 7598 3 7620 1 7618 OAI21X2 $T=1971420 896560 1 0 $X=1971418 $Y=891120
X507 8325 8162 3 8385 1 8401 OAI21X2 $T=2136420 846160 1 180 $X=2131140 $Y=845758
X508 8500 260 3 8502 1 8523 OAI21X2 $T=2152260 967120 1 0 $X=2152258 $Y=961680
X509 8637 260 3 8634 1 8639 OAI21X2 $T=2188560 846160 1 180 $X=2183280 $Y=845758
X510 342 260 3 274 1 275 OAI21X2 $T=2196480 977200 1 180 $X=2191200 $Y=976798
X511 8764 260 3 8782 1 8760 OAI21X2 $T=2206380 846160 0 0 $X=2206378 $Y=845758
X512 8812 260 3 8828 1 8830 OAI21X2 $T=2216940 846160 0 0 $X=2216938 $Y=845758
X513 5286 155 5402 3 1 XNOR2X4 $T=1493580 886480 1 0 $X=1493578 $Y=881040
X514 5831 5835 5901 3 1 XNOR2X4 $T=1591920 785680 0 0 $X=1591918 $Y=785278
X515 5708 6005 6144 3 1 XNOR2X4 $T=1638780 785680 1 0 $X=1638778 $Y=780240
X516 6079 166 6193 3 1 XNOR2X4 $T=1648020 795760 1 0 $X=1648018 $Y=790320
X517 6125 6143 6167 3 1 XNOR2X4 $T=1655940 775600 0 0 $X=1655938 $Y=775198
X518 200 6232 6273 3 1 XNOR2X4 $T=1680360 745360 0 0 $X=1680358 $Y=744958
X519 7315 7335 230 3 1 XNOR2X4 $T=1907400 856240 0 0 $X=1907398 $Y=855838
X520 7452 7473 236 3 1 XNOR2X4 $T=1943700 936880 0 0 $X=1943698 $Y=936478
X521 7676 7574 242 3 1 XNOR2X4 $T=1985940 906640 1 0 $X=1985938 $Y=901200
X522 8545 8523 7977 3 1 XNOR2X4 $T=2162820 957040 1 180 $X=2151600 $Y=956638
X523 8659 8639 7975 3 1 XNOR2X4 $T=2191200 836080 1 180 $X=2179980 $Y=835678
X524 8681 275 7969 3 1 XNOR2X4 $T=2197800 957040 1 180 $X=2186580 $Y=956638
X525 8835 8830 8112 3 1 XNOR2X4 $T=2225520 826000 0 180 $X=2214300 $Y=820560
X526 5538 3 5521 5523 1 5589 OAI21X4 $T=1556280 856240 1 180 $X=1549020 $Y=855838
X527 5673 3 5678 5580 1 5677 OAI21X4 $T=1565520 826000 0 180 $X=1558260 $Y=820560
X528 5729 3 5672 5539 1 5716 OAI21X4 $T=1576740 775600 1 180 $X=1569480 $Y=775198
X529 165 3 5713 5756 1 5731 OAI21X4 $T=1584000 957040 1 180 $X=1576740 $Y=956638
X530 5845 3 166 5895 1 5914 OAI21X4 $T=1597860 765520 1 0 $X=1597858 $Y=760080
X531 5833 3 166 5789 1 5835 OAI21X4 $T=1597860 775600 0 0 $X=1597858 $Y=775198
X532 5649 3 166 5729 1 6005 OAI21X4 $T=1633500 785680 0 180 $X=1626240 $Y=780240
X533 5936 3 166 6158 1 6143 OAI21X4 $T=1657920 765520 0 0 $X=1657918 $Y=765118
X534 166 3 6162 6068 1 6232 OAI21X4 $T=1665180 745360 0 0 $X=1665178 $Y=744958
X535 7082 3 7084 7105 1 7149 OAI21X4 $T=1857900 866320 0 0 $X=1857898 $Y=865918
X536 222 3 7131 7147 1 7080 OAI21X4 $T=1867800 946960 0 0 $X=1867798 $Y=946558
X537 7490 3 7528 7454 1 7473 OAI21X4 $T=1952940 926800 0 180 $X=1945680 $Y=921360
X538 7551 3 7303 7573 1 7577 OAI21X4 $T=1958880 826000 0 0 $X=1958878 $Y=825598
X539 7622 3 7621 7649 1 7712 OAI21X4 $T=1976700 946960 1 0 $X=1976698 $Y=941520
X540 7717 3 7666 7664 1 7480 OAI21X4 $T=1995180 805840 1 180 $X=1987920 $Y=805438
X541 49 3379 1 3 3476 XOR2X2 $T=1135200 856240 1 0 $X=1135198 $Y=850800
X542 3664 97 1 3 3936 XOR2X2 $T=1188000 967120 1 0 $X=1187998 $Y=961680
X543 3382 75 1 3 102 XOR2X2 $T=1200540 946960 0 0 $X=1200538 $Y=946558
X544 117 118 1 3 123 XOR2X2 $T=1336500 977200 1 0 $X=1336498 $Y=971760
X545 119 4561 1 3 125 XOR2X2 $T=1341780 916720 1 0 $X=1341778 $Y=911280
X546 116 115 1 3 143 XOR2X2 $T=1348380 936880 1 0 $X=1348378 $Y=931440
X547 5197 5214 1 3 5430 XOR2X2 $T=1473780 836080 0 0 $X=1473778 $Y=835678
X548 5077 5248 1 3 5364 XOR2X2 $T=1483020 826000 0 0 $X=1483018 $Y=825598
X549 5218 5122 1 3 5267 XOR2X2 $T=1483680 785680 0 0 $X=1483678 $Y=785278
X550 5177 5293 1 3 5401 XOR2X2 $T=1495560 876400 1 0 $X=1495558 $Y=870960
X551 5139 5215 1 3 5410 XOR2X2 $T=1505460 775600 0 0 $X=1505458 $Y=775198
X552 159 5403 1 3 163 XOR2X2 $T=1520640 977200 0 0 $X=1520638 $Y=976798
X553 5544 5685 1 3 5966 XOR2X2 $T=1564200 876400 0 0 $X=1564198 $Y=875998
X554 5759 5755 1 3 5962 XOR2X2 $T=1579380 856240 1 0 $X=1579378 $Y=850800
X555 345 5815 1 3 5965 XOR2X2 $T=1599180 977200 0 0 $X=1599178 $Y=976798
X556 6945 6948 1 3 219 XOR2X2 $T=1833480 946960 1 0 $X=1833478 $Y=941520
X557 7013 6991 1 3 221 XOR2X2 $T=1846680 936880 1 0 $X=1846678 $Y=931440
X558 7214 7258 1 3 228 XOR2X2 $T=1896180 866320 1 0 $X=1896178 $Y=860880
X559 7713 7527 1 3 244 XOR2X2 $T=1993200 836080 0 0 $X=1993198 $Y=835678
X560 7838 7836 1 3 7640 XOR2X2 $T=2016300 906640 1 180 $X=2009700 $Y=906238
X561 247 7877 1 3 6927 XOR2X2 $T=2024880 936880 1 180 $X=2018280 $Y=936478
X562 7908 7904 1 3 6901 XOR2X2 $T=2032140 926800 1 180 $X=2025540 $Y=926398
X563 8200 8162 1 3 8141 XOR2X2 $T=2095500 836080 0 180 $X=2088900 $Y=830640
X564 8390 260 1 3 7901 XOR2X2 $T=2132460 967120 1 180 $X=2125860 $Y=966718
X565 8762 8760 1 3 8266 XOR2X2 $T=2209020 836080 0 180 $X=2202420 $Y=830640
X566 4028 3 4193 1 INVX2 $T=1250700 755440 0 0 $X=1250698 $Y=755038
X567 4496 3 122 1 INVX2 $T=1331880 745360 1 0 $X=1331878 $Y=739920
X568 151 3 5318 1 INVX2 $T=1497540 775600 1 180 $X=1495560 $Y=775198
X569 165 3 5815 1 INVX2 $T=1584660 977200 1 0 $X=1584658 $Y=971760
X570 7149 3 7258 1 INVX2 $T=1898160 856240 1 0 $X=1898158 $Y=850800
X571 7375 3 7427 1 INVX2 $T=1929180 876400 1 180 $X=1927200 $Y=875998
X572 7454 3 7429 1 INVX2 $T=1945680 896560 0 0 $X=1945678 $Y=896158
X573 7480 3 7486 1 INVX2 $T=1950960 805840 0 0 $X=1950958 $Y=805438
X574 7969 3 7967 1 INVX2 $T=2042040 946960 1 0 $X=2042038 $Y=941520
X575 2712 1 3 2713 INVXL $T=953040 946960 1 180 $X=951720 $Y=946558
X576 2820 1 3 2799 INVXL $T=995280 936880 1 180 $X=993960 $Y=936478
X577 77 1 3 3388 INVXL $T=1112760 936880 0 0 $X=1112758 $Y=936478
X578 3319 1 3 3428 INVXL $T=1128600 946960 0 0 $X=1128598 $Y=946558
X579 3381 1 3 3866 INVXL $T=1205820 856240 1 0 $X=1205818 $Y=850800
X580 3963 1 3 4174 INVXL $T=1248720 785680 1 0 $X=1248718 $Y=780240
X581 4306 1 3 4276 INVXL $T=1285680 775600 0 180 $X=1284360 $Y=770160
X582 5497 1 3 5577 INVXL $T=1549680 755440 0 180 $X=1548360 $Y=750000
X583 5538 1 3 5629 INVXL $T=1551000 886480 0 0 $X=1550998 $Y=886078
X584 5516 1 3 5773 INVXL $T=1582020 755440 0 0 $X=1582018 $Y=755038
X585 5716 1 3 5789 INVXL $T=1582020 775600 0 0 $X=1582018 $Y=775198
X586 181 1 3 5943 INVXL $T=1633500 745360 1 180 $X=1632180 $Y=744958
X587 7233 1 3 7231 INVXL $T=1894860 896560 1 180 $X=1893540 $Y=896158
X588 7835 1 3 7809 INVXL $T=2007060 866320 1 180 $X=2005740 $Y=865918
X589 7833 1 3 7855 INVXL $T=2018940 866320 1 0 $X=2018938 $Y=860880
X590 7880 1 3 7927 INVXL $T=2032140 826000 0 0 $X=2032138 $Y=825598
X591 7901 1 3 8048 INVXL $T=2062500 957040 0 180 $X=2061180 $Y=951600
X592 8267 1 3 8269 INVXL $T=2099460 866320 0 180 $X=2098140 $Y=860880
X593 8836 1 3 8856 INVXL $T=2232120 866320 0 180 $X=2230800 $Y=860880
X594 8878 1 3 8829 INVXL $T=2234760 856240 1 180 $X=2233440 $Y=855838
X595 3872 3875 3763 1 3882 3881 3 AOI31X1 $T=1207140 826000 1 0 $X=1207138 $Y=820560
X596 3763 3875 3872 1 3882 3919 3 AOI31X1 $T=1219680 826000 0 180 $X=1216380 $Y=820560
X597 108 4172 4113 1 4130 4170 3 AOI31X1 $T=1254000 916720 1 180 $X=1250700 $Y=916318
X598 224 7177 223 1 7153 7104 3 AOI31X1 $T=1878360 967120 0 0 $X=1878358 $Y=966718
X599 8117 8142 8140 1 8135 7836 3 AOI31X1 $T=2080980 906640 1 180 $X=2077680 $Y=906238
X600 2738 2737 1 3 56 XNOR2X2 $T=966900 957040 1 180 $X=959640 $Y=956638
X601 5179 5360 1 3 5400 XNOR2X2 $T=1499520 795760 0 0 $X=1499518 $Y=795358
X602 5381 5406 1 3 5627 XNOR2X2 $T=1520640 946960 0 0 $X=1520638 $Y=946558
X603 5726 5688 1 3 5963 XNOR2X2 $T=1570800 906640 1 0 $X=1570798 $Y=901200
X604 5775 5731 1 3 5964 XNOR2X2 $T=1582020 946960 1 0 $X=1582018 $Y=941520
X605 5834 5818 1 3 5939 XNOR2X2 $T=1592580 926800 0 0 $X=1592578 $Y=926398
X606 7152 7106 1 3 225 XNOR2X2 $T=1871760 896560 1 0 $X=1871758 $Y=891120
X607 7714 7712 1 3 243 XNOR2X2 $T=1992540 946960 0 0 $X=1992538 $Y=946558
X608 8347 8346 1 3 8003 XNOR2X2 $T=2121900 856240 1 180 $X=2114640 $Y=855838
X609 8412 8401 1 3 8092 XNOR2X2 $T=2138400 826000 1 180 $X=2131140 $Y=825598
X610 8574 8573 1 3 7939 XNOR2X2 $T=2172060 846160 1 180 $X=2164800 $Y=845758
X611 2640 46 3 1 53 XOR2X1 $T=949740 957040 1 180 $X=944460 $Y=956638
X612 2756 2755 3 1 57 XOR2X1 $T=968220 916720 1 180 $X=962940 $Y=916318
X613 3213 75 3 1 3251 XOR2X1 $T=1085700 866320 1 0 $X=1085698 $Y=860880
X614 3343 3342 3 1 3321 XOR2X1 $T=1111440 896560 1 180 $X=1106160 $Y=896158
X615 3034 3379 3 1 3338 XOR2X1 $T=1118700 846160 1 180 $X=1113420 $Y=845758
X616 75 3425 3 1 3391 XOR2X1 $T=1130580 876400 1 180 $X=1125300 $Y=875998
X617 87 86 3 1 3477 XOR2X1 $T=1145100 967120 1 180 $X=1139820 $Y=966718
X618 71 3425 3 1 3665 XOR2X1 $T=1160940 896560 0 0 $X=1160938 $Y=896158
X619 91 74 3 1 3668 XOR2X1 $T=1161600 967120 1 0 $X=1161598 $Y=961680
X620 3885 3644 3 1 3947 XOR2X1 $T=1209780 957040 0 0 $X=1209778 $Y=956638
X621 104 3947 3 1 4080 XOR2X1 $T=1218360 967120 1 0 $X=1218358 $Y=961680
X622 4052 4077 3 1 3848 XOR2X1 $T=1241460 775600 1 180 $X=1236180 $Y=775198
X623 3963 4082 3 1 4052 XOR2X1 $T=1242780 785680 1 180 $X=1237500 $Y=785278
X624 65 3035 3 1 110 XOR2X1 $T=1240140 805840 0 0 $X=1240138 $Y=805438
X625 4082 63 3 1 4244 XOR2X1 $T=1265220 886480 1 0 $X=1265218 $Y=881040
X626 4188 4218 3 1 4413 XOR2X1 $T=1272480 745360 1 0 $X=1272478 $Y=739920
X627 4261 108 3 1 4274 XOR2X1 $T=1273140 977200 1 0 $X=1273138 $Y=971760
X628 4328 4307 3 1 4359 XOR2X1 $T=1290960 866320 0 0 $X=1290958 $Y=865918
X629 4346 4300 3 1 112 XOR2X1 $T=1292280 785680 0 0 $X=1292278 $Y=785278
X630 5008 5118 3 1 159 XOR2X1 $T=1479720 977200 1 0 $X=1479718 $Y=971760
X631 5072 5282 3 1 5381 XOR2X1 $T=1490280 946960 0 0 $X=1490278 $Y=946558
X632 5071 5362 3 1 5429 XOR2X1 $T=1504140 745360 0 0 $X=1504138 $Y=744958
X633 5279 5405 3 1 5547 XOR2X1 $T=1511400 936880 1 0 $X=1511398 $Y=931440
X634 7103 7104 3 1 220 XOR2X1 $T=1863180 977200 0 180 $X=1857900 $Y=971760
X635 7834 7810 3 1 7234 XOR2X1 $T=2013000 957040 1 180 $X=2007720 $Y=956638
X636 7835 7833 3 1 7446 XOR2X1 $T=2013660 866320 0 180 $X=2008380 $Y=860880
X637 7975 7941 3 1 7317 XOR2X1 $T=2045340 815920 0 180 $X=2040060 $Y=810480
X638 346 248 3 1 7834 XOR2X1 $T=2047980 977200 1 180 $X=2042700 $Y=976798
X639 2798 1 2797 2756 3 NOR2BX1 $T=978780 916720 1 180 $X=976140 $Y=916318
X640 3460 1 3478 3462 3 NOR2BX1 $T=1137180 916720 0 0 $X=1137178 $Y=916318
X641 5219 1 5125 5239 3 NOR2BX1 $T=1479720 826000 1 0 $X=1479718 $Y=820560
X642 153 1 152 5260 3 NOR2BX1 $T=1485000 745360 0 0 $X=1484998 $Y=744958
X643 5379 1 5315 5407 3 NOR2BX1 $T=1506780 936880 0 0 $X=1506778 $Y=936478
X644 5590 1 5455 5709 3 NOR2BX1 $T=1566180 836080 1 0 $X=1566178 $Y=830640
X645 5729 1 5649 6079 3 NOR2BX1 $T=1631520 795760 1 0 $X=1631518 $Y=790320
X646 182 1 174 6069 3 NOR2BX1 $T=1634820 745360 1 0 $X=1634818 $Y=739920
X647 6900 1 6898 6945 3 NOR2BX1 $T=1831500 916720 0 0 $X=1831498 $Y=916318
X648 7494 1 7388 7489 3 NOR2BX1 $T=1951620 815920 1 180 $X=1948980 $Y=815518
X649 7717 1 7644 7713 3 NOR2BX1 $T=1995840 815920 1 180 $X=1993200 $Y=815518
X650 8746 1 8758 8761 3 NOR2BX1 $T=2204400 866320 1 0 $X=2204398 $Y=860880
X651 8741 1 8743 8762 3 NOR2BX1 $T=2208360 886480 1 180 $X=2205720 $Y=886078
X652 8657 1 8758 8766 3 NOR2BX1 $T=2212320 866320 1 180 $X=2209680 $Y=865918
X653 63 62 2946 2615 1 3 2841 ADDFX2 $T=1017720 916720 0 180 $X=1003860 $Y=911280
X654 3033 3035 3016 2825 1 3 2865 ADDFX2 $T=1036860 906640 0 180 $X=1023000 $Y=901200
X655 3127 3072 3053 2886 1 3 64 ADDFX2 $T=1049400 957040 1 180 $X=1035540 $Y=956638
X656 3190 3135 3128 2864 1 3 2884 ADDFX2 $T=1059960 936880 0 180 $X=1046100 $Y=931440
X657 71 65 3155 2505 1 3 2695 ADDFX2 $T=1070520 916720 0 180 $X=1056660 $Y=911280
X658 70 69 3156 3053 1 3 67 ADDFX2 $T=1073160 967120 0 180 $X=1059300 $Y=961680
X659 72 3035 3157 3128 1 3 3127 ADDFX2 $T=1074480 926800 1 180 $X=1060620 $Y=926398
X660 79 62 68 3072 1 3 66 ADDFX2 $T=1075800 977200 0 180 $X=1061940 $Y=971760
X661 3155 75 69 3016 1 3 3190 ADDFX2 $T=1090320 906640 1 180 $X=1076460 $Y=906238
X662 72 65 76 3156 1 3 73 ADDFX2 $T=1096920 967120 0 180 $X=1083060 $Y=961680
X663 124 126 133 4716 1 3 129 ADDFX2 $T=1357620 977200 0 0 $X=1357618 $Y=976798
X664 127 131 135 4770 1 3 141 ADDFX2 $T=1373460 967120 0 0 $X=1373458 $Y=966718
X665 130 4752 4770 4791 1 3 4771 ADDFX2 $T=1375440 936880 0 0 $X=1375438 $Y=936478
X666 4751 134 4790 4795 1 3 4817 ADDFX2 $T=1378080 876400 1 0 $X=1378078 $Y=870960
X667 133 139 138 4768 1 3 4752 ADDFX2 $T=1393920 926800 1 180 $X=1380060 $Y=926398
X668 133 138 136 4813 1 3 4790 ADDFX2 $T=1381380 866320 1 0 $X=1381378 $Y=860880
X669 136 128 130 4814 1 3 4789 ADDFX2 $T=1382700 815920 1 0 $X=1382698 $Y=810480
X670 135 137 123 4816 1 3 4792 ADDFX2 $T=1383360 836080 0 0 $X=1383358 $Y=835678
X671 4789 143 4816 4835 1 3 4885 ADDFX2 $T=1386660 826000 1 0 $X=1386658 $Y=820560
X672 4792 125 4795 4836 1 3 4886 ADDFX2 $T=1387320 846160 0 0 $X=1387318 $Y=845758
X673 4767 132 4904 4909 1 3 4948 ADDFX2 $T=1397880 896560 0 0 $X=1397878 $Y=896158
X674 4835 4889 4906 4921 1 3 4944 ADDFX2 $T=1398540 795760 0 0 $X=1398538 $Y=795358
X675 4814 120 125 4907 1 3 4906 ADDFX2 $T=1399200 785680 0 0 $X=1399198 $Y=785278
X676 4884 4891 4907 4923 1 3 4981 ADDFX2 $T=1399860 785680 1 0 $X=1399858 $Y=780240
X677 136 4768 4837 4904 1 3 4970 ADDFX2 $T=1399860 916720 1 0 $X=1399858 $Y=911280
X678 128 4716 136 4924 1 3 4930 ADDFX2 $T=1400520 957040 1 0 $X=1400518 $Y=951600
X679 4887 143 4817 4925 1 3 5054 ADDFX2 $T=1401180 876400 1 0 $X=1401178 $Y=870960
X680 132 135 143 4890 1 3 4884 ADDFX2 $T=1415040 765520 1 180 $X=1401180 $Y=765118
X681 134 133 123 4891 1 3 4889 ADDFX2 $T=1416360 815920 1 180 $X=1402500 $Y=815518
X682 132 143 120 146 1 3 4984 ADDFX2 $T=1404480 745360 1 0 $X=1404478 $Y=739920
X683 143 134 4791 4949 1 3 5057 ADDFX2 $T=1407780 936880 1 0 $X=1407778 $Y=931440
X684 132 4813 120 4922 1 3 4901 ADDFX2 $T=1421640 866320 0 180 $X=1407780 $Y=860880
X685 4905 125 4890 4958 1 3 4966 ADDFX2 $T=1409760 775600 1 0 $X=1409758 $Y=770160
X686 130 136 120 4959 1 3 4905 ADDFX2 $T=1409760 805840 0 0 $X=1409758 $Y=805438
X687 4885 4922 4836 4947 1 3 5023 ADDFX2 $T=1410420 836080 0 0 $X=1410418 $Y=835678
X688 4930 123 147 4983 1 3 5004 ADDFX2 $T=1415040 967120 1 0 $X=1415038 $Y=961680
X689 123 134 4959 4987 1 3 5038 ADDFX2 $T=1418340 805840 1 0 $X=1418338 $Y=800400
X690 5010 4983 4903 5072 1 3 5118 ADDFX2 $T=1436160 957040 1 0 $X=1436158 $Y=951600
X691 8282 258 8348 8264 1 3 8326 ADDFX2 $T=2129820 916720 0 180 $X=2115960 $Y=911280
X692 8519 8282 8394 8328 1 3 8389 ADDFX2 $T=2144340 896560 1 180 $X=2130480 $Y=896158
X693 257 263 261 8348 1 3 8394 ADDFX2 $T=2145000 926800 1 180 $X=2131140 $Y=926398
X694 8522 8501 8467 8443 1 3 8445 ADDFX2 $T=2158860 916720 1 180 $X=2145000 $Y=916318
X695 258 267 259 8501 1 3 8550 ADDFX2 $T=2151600 946960 1 0 $X=2151598 $Y=941520
X696 269 261 8550 8467 1 3 8742 ADDFX2 $T=2156220 926800 1 0 $X=2156218 $Y=921360
X697 276 265 261 8763 1 3 8759 ADDFX2 $T=2197140 926800 0 0 $X=2197138 $Y=926398
X698 8793 8763 8742 8462 1 3 8698 ADDFX2 $T=2211000 916720 0 180 $X=2197140 $Y=911280
X699 8744 8759 8784 8791 1 3 8792 ADDFX2 $T=2201760 916720 0 0 $X=2201758 $Y=916318
X700 276 265 257 8788 1 3 8805 ADDFX2 $T=2203080 957040 1 0 $X=2203078 $Y=951600
X701 272 277 8788 8793 1 3 8784 ADDFX2 $T=2203740 946960 1 0 $X=2203738 $Y=941520
X702 284 283 8875 8860 1 3 8810 ADDFX2 $T=2242020 967120 1 180 $X=2228160 $Y=966718
X703 272 280 8861 8900 1 3 8875 ADDFX2 $T=2228820 957040 1 0 $X=2228818 $Y=951600
X704 279 281 8896 8895 1 3 8915 ADDFX2 $T=2228820 967120 1 0 $X=2228818 $Y=961680
X705 285 269 8877 8744 1 3 8857 ADDFX2 $T=2242680 936880 0 180 $X=2228820 $Y=931440
X706 2504 2505 3 1 2565 XNOR2X1 $T=920040 957040 0 0 $X=920038 $Y=956638
X707 2547 2548 3 1 51 XNOR2X1 $T=933240 926800 1 180 $X=927960 $Y=926398
X708 2565 2567 3 1 52 XNOR2X1 $T=933240 957040 0 0 $X=933238 $Y=956638
X709 71 3155 3 1 3213 XNOR2X1 $T=1073160 866320 1 0 $X=1073158 $Y=860880
X710 3251 3485 3 1 3619 XNOR2X1 $T=1139820 795760 1 0 $X=1139818 $Y=790320
X711 49 63 3 1 3482 XNOR2X1 $T=1147740 926800 1 180 $X=1142460 $Y=926398
X712 110 3034 3 1 4077 XNOR2X1 $T=1258620 805840 0 180 $X=1253340 $Y=800400
X713 4138 4187 3 1 4333 XNOR2X1 $T=1254660 896560 0 0 $X=1254658 $Y=896158
X714 4082 65 3 1 4346 XNOR2X1 $T=1283700 805840 1 0 $X=1283698 $Y=800400
X715 5055 5116 3 1 5177 XNOR2X1 $T=1454640 866320 0 0 $X=1454638 $Y=865918
X716 5163 5220 3 1 5279 XNOR2X1 $T=1479720 936880 1 0 $X=1479718 $Y=931440
X717 8113 8110 3 1 7924 XNOR2X1 $T=2074380 896560 0 180 $X=2069100 $Y=891120
X718 8121 8120 3 1 7996 XNOR2X1 $T=2076360 876400 1 180 $X=2071080 $Y=875998
X719 5155 151 3 5134 1 4994 5039 5159 OAI221XL $T=1466520 785680 1 180 $X=1461900 $Y=785278
X720 50 2504 49 1 3 43 ADDHXL $T=925980 967120 1 180 $X=918720 $Y=966718
X721 50 3033 3034 1 3 2946 ADDHXL $T=1026300 916720 1 0 $X=1026298 $Y=911280
X722 74 3157 65 1 3 3135 ADDHXL $T=1087020 926800 1 180 $X=1079760 $Y=926398
X723 185 6046 188 1 3 6090 ADDHXL $T=1636800 957040 0 0 $X=1636798 $Y=956638
X724 6090 6118 183 1 3 6152 ADDHXL $T=1649340 957040 0 0 $X=1649338 $Y=956638
X725 6156 6160 190 1 3 6168 ADDHXL $T=1659240 946960 0 0 $X=1659238 $Y=946558
X726 6152 196 194 1 3 6156 ADDHXL $T=1669140 957040 1 180 $X=1661880 $Y=956638
X727 6168 6185 184 1 3 6205 ADDHXL $T=1663200 936880 0 0 $X=1663198 $Y=936478
X728 6205 6208 199 1 3 6291 ADDHXL $T=1681680 936880 0 0 $X=1681678 $Y=936478
X729 6291 6316 202 1 3 6370 ADDHXL $T=1694220 936880 0 0 $X=1694218 $Y=936478
X730 6301 6369 210 1 3 211 ADDHXL $T=1696860 967120 0 0 $X=1696858 $Y=966718
X731 6370 6368 203 1 3 6301 ADDHXL $T=1704120 946960 1 180 $X=1696860 $Y=946558
X732 1 42 43 44 3 NOR2XL $T=894300 977200 0 0 $X=894298 $Y=976798
X733 1 4082 72 4307 3 NOR2XL $T=1278420 866320 0 0 $X=1278418 $Y=865918
X734 1 5155 152 5200 3 NOR2XL $T=1469160 785680 0 0 $X=1469158 $Y=785278
X735 1 8218 255 8179 3 NOR2XL $T=2096820 926800 1 180 $X=2094840 $Y=926398
X736 1 8325 8324 8305 3 NOR2XL $T=2117280 866320 1 180 $X=2115300 $Y=865918
X737 3319 77 3359 3 1 3320 XOR3X2 $T=1101540 946960 0 0 $X=1101538 $Y=946558
X738 82 3035 75 3 1 3343 XOR3X2 $T=1127940 916720 0 180 $X=1116060 $Y=911280
X739 3341 3345 3321 3 1 3424 XOR3X2 $T=1117380 826000 0 0 $X=1117378 $Y=825598
X740 85 3476 3477 3 1 3573 XOR3X2 $T=1142460 866320 0 0 $X=1142458 $Y=865918
X741 93 3483 3668 3 1 3664 XOR3X2 $T=1184040 957040 1 180 $X=1172160 $Y=956638
X742 3661 3724 3339 3 1 3746 XOR3X2 $T=1178100 815920 0 0 $X=1178098 $Y=815518
X743 3520 3787 3573 3 1 3915 XOR3X2 $T=1192620 886480 1 0 $X=1192618 $Y=881040
X744 99 3665 100 3 1 3867 XOR3X2 $T=1192620 936880 0 0 $X=1192618 $Y=936478
X745 3872 3844 3801 3 1 3980 XOR3X2 $T=1213740 866320 1 0 $X=1213738 $Y=860880
X746 3725 3381 4071 3 1 4085 XOR3X2 $T=1228920 846160 0 0 $X=1228918 $Y=845758
X747 89 4233 4244 3 1 4194 XOR3X2 $T=1259940 815920 0 0 $X=1259938 $Y=815518
X748 8270 8264 8207 3 1 7835 XOR3X2 $T=2106720 866320 1 180 $X=2094840 $Y=865918
X749 77 3319 1 3359 3 3389 AOI21XL $T=1120020 946960 0 0 $X=1120018 $Y=946558
X750 3503 3479 1 3506 3 3571 AOI21XL $T=1143780 775600 0 0 $X=1143778 $Y=775198
X751 3345 3321 3341 3 3337 1 OAI2BB1X1 $T=1112100 836080 0 180 $X=1108800 $Y=830640
X752 3338 3320 3346 3 3340 1 OAI2BB1X1 $T=1112760 866320 0 180 $X=1109460 $Y=860880
X753 3382 3391 3383 3 3362 1 OAI2BB1X1 $T=1120020 876400 1 180 $X=1116720 $Y=875998
X754 80 3343 72 3 3406 1 OAI2BB1X1 $T=1124640 906640 1 0 $X=1124638 $Y=901200
X755 83 82 81 3 3383 1 OAI2BB1X1 $T=1127940 926800 0 180 $X=1124640 $Y=921360
X756 3455 3251 3452 3 3446 1 OAI2BB1X1 $T=1135860 805840 0 180 $X=1132560 $Y=800400
X757 3476 3477 85 3 3456 1 OAI2BB1X1 $T=1142460 856240 1 180 $X=1139160 $Y=855838
X758 3572 3457 3570 3 3592 1 OAI2BB1X1 $T=1153020 846160 1 0 $X=1153018 $Y=840720
X759 78 63 76 3 3594 1 OAI2BB1X1 $T=1156320 957040 1 0 $X=1156318 $Y=951600
X760 3425 3034 69 3 3641 1 OAI2BB1X1 $T=1162920 886480 1 0 $X=1162918 $Y=881040
X761 86 76 3642 3 3645 1 OAI2BB1X1 $T=1164240 926800 1 0 $X=1164238 $Y=921360
X762 3670 3687 3645 3 3692 1 OAI2BB1X1 $T=1174800 876400 0 0 $X=1174798 $Y=875998
X763 3689 3668 93 3 3693 1 OAI2BB1X1 $T=1177440 946960 0 0 $X=1177438 $Y=946558
X764 96 3664 95 3 3704 1 OAI2BB1X1 $T=1183380 977200 0 180 $X=1180080 $Y=971760
X765 100 3665 99 3 3789 1 OAI2BB1X1 $T=1195260 926800 0 0 $X=1195258 $Y=926398
X766 3573 3787 3785 3 3801 1 OAI2BB1X1 $T=1196580 866320 0 0 $X=1196578 $Y=865918
X767 3867 3845 3838 3 3908 1 OAI2BB1X1 $T=1208460 916720 0 0 $X=1208458 $Y=916318
X768 3967 104 3644 3 4006 1 OAI2BB1X1 $T=1221660 957040 1 0 $X=1221658 $Y=951600
X769 4233 4244 89 3 4298 1 OAI2BB1X1 $T=1279080 826000 1 0 $X=1279078 $Y=820560
X770 71 4307 4345 3 111 1 OAI2BB1X1 $T=1292280 866320 1 0 $X=1292278 $Y=860880
X771 5137 5160 5029 3 5222 1 OAI2BB1X1 $T=1462560 826000 1 0 $X=1462558 $Y=820560
X772 5760 5731 5680 3 5818 1 OAI2BB1X1 $T=1580040 926800 0 0 $X=1580038 $Y=926398
X773 178 170 6002 3 6023 1 OAI2BB1X1 $T=1629540 856240 1 0 $X=1629538 $Y=850800
X774 178 172 6003 3 6037 1 OAI2BB1X1 $T=1629540 866320 0 0 $X=1629538 $Y=865918
X775 178 167 6027 3 6039 1 OAI2BB1X1 $T=1634820 886480 1 0 $X=1634818 $Y=881040
X776 178 177 6076 3 5999 1 OAI2BB1X1 $T=1648680 846160 0 180 $X=1645380 $Y=840720
X777 178 187 6142 3 6048 1 OAI2BB1X1 $T=1659240 846160 0 180 $X=1655940 $Y=840720
X778 178 186 6159 3 6268 1 OAI2BB1X1 $T=1661220 876400 0 0 $X=1661218 $Y=875998
X779 178 197 6204 3 6155 1 OAI2BB1X1 $T=1675080 846160 0 180 $X=1671780 $Y=840720
X780 178 206 6249 3 6243 1 OAI2BB1X1 $T=1687620 846160 0 180 $X=1684320 $Y=840720
X781 178 213 6373 3 6372 1 OAI2BB1X1 $T=1706100 846160 0 180 $X=1702800 $Y=840720
X782 178 216 6428 3 6443 1 OAI2BB1X1 $T=1718640 856240 1 0 $X=1718638 $Y=850800
X783 178 215 6404 3 6442 1 OAI2BB1X1 $T=1718640 866320 1 0 $X=1718638 $Y=860880
X784 178 214 6429 3 6425 1 OAI2BB1X1 $T=1718640 886480 1 0 $X=1718638 $Y=881040
X785 246 245 7810 3 7238 1 OAI2BB1X1 $T=2009700 977200 1 180 $X=2006400 $Y=976798
X786 7896 7924 7907 3 7637 1 OAI2BB1X1 $T=2032140 886480 0 180 $X=2028840 $Y=881040
X787 7941 7975 8111 3 7978 1 OAI2BB1X1 $T=2075040 815920 1 180 $X=2071740 $Y=815518
X788 8117 8139 8122 3 8135 1 OAI2BB1X1 $T=2086920 906640 1 180 $X=2083620 $Y=906238
X789 8850 8638 8746 3 8786 1 OAI2BB1X1 $T=2228160 866320 0 180 $X=2224860 $Y=860880
X790 2820 3 2800 1 2738 NAND2BXL $T=981420 936880 1 180 $X=978780 $Y=936478
X791 3849 3 3617 1 3904 NAND2BXL $T=1210440 765520 0 0 $X=1210438 $Y=765118
X792 4213 3 4222 1 4218 NAND2BXL $T=1267860 745360 0 180 $X=1265220 $Y=739920
X793 4957 3 5022 1 5077 NAND2BXL $T=1445400 826000 1 0 $X=1445398 $Y=820560
X794 5513 3 5452 1 5628 NAND2BXL $T=1538460 815920 0 0 $X=1538458 $Y=815518
X795 5679 3 5674 1 5834 NAND2BXL $T=1564200 906640 0 0 $X=1564198 $Y=906238
X796 8146 3 8092 1 8090 NAND2BXL $T=2082300 805840 1 180 $X=2079660 $Y=805438
X797 272 8282 3 1 CLKBUFX3 $T=2184600 936880 0 180 $X=2181960 $Y=931440
X798 44 2397 42 43 1 3 48 AOI2BB2X1 $T=899580 977200 0 0 $X=899578 $Y=976798
X799 49 89 3034 4240 1 3 4233 AOI2BB2X1 $T=1266540 826000 0 0 $X=1266538 $Y=825598
X800 127 128 130 4751 1 3 4767 ADDFHX1 $T=1365540 896560 0 0 $X=1365538 $Y=896158
X801 126 137 135 4793 1 3 4837 ADDFHX1 $T=1375440 916720 1 0 $X=1375438 $Y=911280
X802 132 4771 4796 4812 1 3 4903 ADDFHX1 $T=1377420 946960 0 0 $X=1377418 $Y=946558
X803 123 4924 143 4988 1 3 5010 ADDFHX1 $T=1414380 936880 0 0 $X=1414378 $Y=936478
X804 4970 125 4988 5035 1 3 5162 ADDFHX1 $T=1425600 916720 1 0 $X=1425598 $Y=911280
X805 8805 8895 8857 8851 1 3 8859 ADDFHX1 $T=2245320 896560 1 180 $X=2230140 $Y=896158
X806 282 8915 8900 8914 1 3 8943 ADDFHX1 $T=2233440 926800 1 0 $X=2233438 $Y=921360
X807 140 3 142 1 4811 4796 NAND3X1 $T=1389300 977200 0 0 $X=1389298 $Y=976798
X808 7997 3 8048 1 7967 8051 NAND3X1 $T=2056560 946960 1 0 $X=2056558 $Y=941520
X809 259 258 257 8218 3 1 8207 CMPR32X1 $T=2111340 936880 1 180 $X=2097480 $Y=936478
X810 263 265 257 8519 3 1 8522 CMPR32X1 $T=2145000 936880 1 0 $X=2144998 $Y=931440
X811 277 259 269 8877 3 1 8896 CMPR32X1 $T=2228820 946960 0 0 $X=2228818 $Y=946558
X812 257 265 272 8861 3 1 347 CMPR32X1 $T=2242680 977200 1 180 $X=2228820 $Y=976798
X813 4793 123 120 4887 1 3 5020 ADDFHX2 $T=1397880 896560 1 0 $X=1397878 $Y=891120
X814 4901 4925 4886 4968 1 3 5116 ADDFHX2 $T=1404480 856240 1 0 $X=1404478 $Y=850800
X815 145 348 5004 5008 1 3 5203 ADDFHX2 $T=1413060 977200 0 0 $X=1413058 $Y=976798
X816 125 5020 4949 5024 1 3 5202 ADDFHX2 $T=1422960 896560 0 0 $X=1422958 $Y=896158
X817 4909 5024 5054 5055 1 3 5123 ADDFHX2 $T=1423620 866320 0 0 $X=1423618 $Y=865918
X818 5057 4812 5162 5163 1 3 5282 ADDFHX2 $T=1444080 926800 0 0 $X=1444078 $Y=926398
X819 4948 5035 5202 5175 1 3 5220 ADDFHX2 $T=1455960 906640 1 0 $X=1455958 $Y=901200
X820 4306 3155 3 1 4285 OR2X1 $T=1283700 775600 1 180 $X=1281060 $Y=775198
X821 188 183 3 1 349 OR2X1 $T=1644720 977200 1 180 $X=1642080 $Y=976798
X822 49 1 3035 3 CLKINVX3 $T=1090980 926800 0 0 $X=1090978 $Y=926398
X823 4038 1 4010 3 CLKINVX3 $T=1244760 876400 0 0 $X=1244758 $Y=875998
X824 3746 1 4452 3 CLKINVX3 $T=1301520 815920 0 0 $X=1301518 $Y=815518
X825 4278 1 4453 3 CLKINVX3 $T=1308120 946960 0 0 $X=1308118 $Y=946558
X826 4413 1 4494 3 CLKINVX3 $T=1324620 745360 1 0 $X=1324618 $Y=739920
X827 164 1 5768 3 CLKINVX3 $T=1568820 977200 1 0 $X=1568818 $Y=971760
X828 181 1 6158 3 CLKINVX3 $T=1668480 755440 0 0 $X=1668478 $Y=755038
X829 7151 1 7175 3 CLKINVX3 $T=1871100 876400 1 180 $X=1869120 $Y=875998
X830 7428 1 7482 3 CLKINVX3 $T=1940400 876400 0 0 $X=1940398 $Y=875998
X831 8004 1 7971 3 CLKINVX3 $T=2046660 815920 1 180 $X=2044680 $Y=815518
X832 8593 1 8640 3 CLKINVX3 $T=2193840 866320 1 0 $X=2193838 $Y=860880
X833 4132 4113 1 4110 3936 4105 3 AOI22X1 $T=1246740 946960 1 180 $X=1243440 $Y=946558
X834 183 6066 1 6050 194 6076 3 AOI22X1 $T=1653960 896560 0 180 $X=1650660 $Y=891120
X835 212 6066 1 6050 207 6404 3 AOI22X1 $T=1710720 906640 0 0 $X=1710718 $Y=906238
X836 8207 8264 1 8267 8268 8178 3 AOI22X1 $T=2100120 876400 0 0 $X=2100118 $Y=875998
X837 8387 8388 1 8326 8328 8370 3 AOI22X1 $T=2132460 886480 1 180 $X=2129160 $Y=886078
X838 3155 4324 4306 4082 3 1 4300 OAI2BB2X1 $T=1288320 785680 1 180 $X=1283700 $Y=785278
X839 3475 3452 3 1 3485 XNOR2XL $T=1141800 805840 1 0 $X=1141798 $Y=800400
X840 3623 3622 3 1 3717 XNOR2XL $T=1162920 785680 0 0 $X=1162918 $Y=785278
X841 3847 3904 3 1 4042 XNOR2XL $T=1210440 775600 0 0 $X=1210438 $Y=775198
X842 3841 3865 3 1 4122 XNOR2XL $T=1219680 795760 1 0 $X=1219678 $Y=790320
X843 71 89 3 1 4328 XNOR2XL $T=1296240 876400 1 180 $X=1290960 $Y=875998
X844 4561 119 120 1 3 OR2X4 $T=1341780 916720 0 0 $X=1341778 $Y=916318
X845 163 4476 5548 1 3 OR2X4 $T=1543080 977200 0 0 $X=1543078 $Y=976798
X846 5961 120 6668 1 3 OR2X4 $T=1772100 906640 0 0 $X=1772098 $Y=906238
X847 5962 7148 7083 1 3 OR2X4 $T=1873740 856240 1 180 $X=1869780 $Y=855838
X848 5966 7150 7085 1 3 OR2X4 $T=1873740 886480 1 180 $X=1869780 $Y=886078
X849 7901 7979 7877 1 3 OR2X4 $T=2046660 957040 0 180 $X=2042700 $Y=951600
X850 7926 8004 7948 1 3 OR2X4 $T=2055900 815920 0 0 $X=2055898 $Y=815518
X851 7969 7968 8049 1 3 OR2X4 $T=2055900 916720 0 0 $X=2055898 $Y=916318
X852 5677 166 3 1 INVX8 $T=1621620 795760 1 0 $X=1621618 $Y=790320
X853 7303 7527 3 1 INVX8 $T=1958880 836080 0 0 $X=1958878 $Y=835678
X854 7577 7528 3 1 INVX8 $T=1965480 906640 0 180 $X=1961520 $Y=901200
X855 7598 7620 7676 3 1 NAND2BX2 $T=1981980 896560 1 0 $X=1981978 $Y=891120
X856 7880 7939 7881 3 1 NAND2BX2 $T=2034780 856240 1 0 $X=2034778 $Y=850800
X857 3764 3841 3743 3847 1 3 OAI2BB1X2 $T=1200540 785680 1 0 $X=1200538 $Y=780240
X858 108 4063 4010 3872 1 3 OAI2BB1X2 $T=1240140 866320 1 180 $X=1235520 $Y=865918
X859 161 160 157 5403 1 3 OAI2BB1X2 $T=1516020 977200 1 180 $X=1511400 $Y=976798
X860 7833 7835 7853 7896 1 3 OAI2BB1X2 $T=2026860 866320 0 0 $X=2026858 $Y=865918
X861 7877 7968 7967 7880 1 3 OAI2BB1X2 $T=2044680 916720 1 180 $X=2040060 $Y=916318
X862 8037 8003 7833 7553 1 3 OAI2BB1X2 $T=2051940 846160 0 180 $X=2047320 $Y=840720
X863 4051 4076 3951 3 1 4188 AND3X2 $T=1239480 765520 0 0 $X=1239478 $Y=765118
X864 4107 4172 4113 3 1 4139 AND3X2 $T=1256640 916720 0 0 $X=1256638 $Y=916318
X865 7978 7948 7976 3 1 7643 AND3X2 $T=2042040 815920 1 180 $X=2038740 $Y=815518
X866 74 89 3461 3 1 NOR2BX2 $T=1154340 826000 1 180 $X=1150380 $Y=825598
X867 247 7904 7968 3 1 NOR2BX2 $T=2052600 926800 1 0 $X=2052598 $Y=921360
X868 80 63 3 1 3342 XOR2XL $T=1121340 896560 1 180 $X=1116060 $Y=896158
X869 3506 3503 3 1 3622 XOR2XL $T=1155000 785680 1 0 $X=1154998 $Y=780240
X870 3665 3034 3 1 3687 XOR2XL $T=1172160 906640 1 0 $X=1172158 $Y=901200
X871 3919 3918 3 1 3952 XOR2XL $T=1215720 815920 0 0 $X=1215718 $Y=815518
X872 1 4169 3998 108 4139 3 NAND3X2 $T=1252680 866320 0 0 $X=1252678 $Y=865918
X873 1 4262 113 4418 4285 3 NAND3X2 $T=1304820 775600 0 0 $X=1304818 $Y=775198
X874 1 8090 7410 8056 8037 3 NAND3X2 $T=2057880 805840 0 0 $X=2057878 $Y=805438
X875 1 8050 8037 8057 7948 3 NAND3X2 $T=2057880 836080 1 0 $X=2057878 $Y=830640
X876 180 179 170 5999 173 1 3 5958 SDFFRHQXL $T=1633500 836080 1 180 $X=1617000 $Y=835678
X877 180 179 172 6023 173 1 3 5944 SDFFRHQXL $T=1639440 846160 0 180 $X=1622940 $Y=840720
X878 180 179 167 6037 173 1 3 5960 SDFFRHQXL $T=1643400 856240 1 180 $X=1626900 $Y=855838
X879 180 179 186 6039 173 1 3 5900 SDFFRHQXL $T=1644060 876400 1 180 $X=1627560 $Y=875998
X880 180 179 190 6077 173 1 3 183 SDFFRHQXL $T=1651320 936880 1 180 $X=1634820 $Y=936478
X881 180 179 177 6048 173 1 3 6120 SDFFRHQXL $T=1637460 836080 0 0 $X=1637458 $Y=835678
X882 180 179 187 6155 173 1 3 6206 SDFFRHQXL $T=1657920 836080 0 0 $X=1657918 $Y=835678
X883 180 179 199 6268 173 1 3 6119 SDFFRHQXL $T=1692240 876400 0 180 $X=1675740 $Y=870960
X884 180 179 197 6243 173 1 3 6290 SDFFRHQXL $T=1677720 836080 0 0 $X=1677718 $Y=835678
X885 180 179 206 6372 173 1 3 6406 SDFFRHQXL $T=1698180 836080 0 0 $X=1698178 $Y=835678
X886 180 179 215 6425 173 1 3 6477 SDFFRHQXL $T=1714680 866320 0 0 $X=1714678 $Y=865918
X887 180 179 216 6442 173 1 3 6481 SDFFRHQXL $T=1716660 846160 1 0 $X=1716658 $Y=840720
X888 180 179 213 6443 173 1 3 6482 SDFFRHQXL $T=1717980 836080 0 0 $X=1717978 $Y=835678
X889 83 1 3034 3 BUFX3 $T=1111440 916720 1 180 $X=1108800 $Y=916318
X890 62 1 4082 3 BUFX3 $T=1269840 896560 1 0 $X=1269838 $Y=891120
X891 5900 1 167 3 BUFX3 $T=1605120 876400 1 180 $X=1602480 $Y=875998
X892 5944 1 170 3 BUFX3 $T=1616340 846160 0 180 $X=1613700 $Y=840720
X893 5960 1 172 3 BUFX3 $T=1618980 856240 1 180 $X=1616340 $Y=855838
X894 5958 1 177 3 BUFX3 $T=1622940 826000 0 0 $X=1622938 $Y=825598
X895 6120 1 187 3 BUFX3 $T=1650660 826000 1 180 $X=1648020 $Y=825598
X896 6119 1 186 3 BUFX3 $T=1653300 866320 0 180 $X=1650660 $Y=860880
X897 6206 1 197 3 BUFX3 $T=1669140 826000 1 180 $X=1666500 $Y=825598
X898 6290 1 206 3 BUFX3 $T=1693560 826000 1 180 $X=1690920 $Y=825598
X899 6482 1 216 3 BUFX3 $T=1733160 826000 0 0 $X=1733158 $Y=825598
X900 6477 1 214 3 BUFX3 $T=1750980 866320 0 0 $X=1750978 $Y=865918
X901 6481 1 215 3 BUFX3 $T=1752300 846160 1 0 $X=1752298 $Y=840720
X902 7876 1 7102 3 BUFX3 $T=2022240 957040 1 0 $X=2022238 $Y=951600
X903 4107 4130 4139 1 108 3 4033 4138 AOI221X1 $T=1252020 906640 0 180 $X=1247400 $Y=901200
X904 110 4415 1 4344 4232 111 110 4306 3 AOI222X2 $T=1295580 745360 1 180 $X=1286340 $Y=744958
X905 4172 1 4132 4261 3 NOR2BXL $T=1275780 967120 1 0 $X=1275778 $Y=961680
X906 3379 1 3623 3619 3 3571 3849 AOI211X1 $T=1169520 775600 0 0 $X=1169518 $Y=775198
X907 75 84 3 1 3449 3359 AOI2BB1X1 $T=1138500 946960 1 180 $X=1135200 $Y=946558
X908 110 111 3 1 4438 4344 AOI2BB1X1 $T=1309440 745360 0 0 $X=1309438 $Y=744958
X909 3449 3482 3479 3462 3 1 MXI2X1 $T=1141800 936880 0 180 $X=1137180 $Y=931440
X910 4049 4053 3 4046 1 4032 4038 OAI211X1 $T=1238820 886480 1 180 $X=1234860 $Y=886078
X911 3320 3346 3338 3 1 3381 XNOR3X2 $T=1106160 856240 1 0 $X=1106158 $Y=850800
X912 3391 3382 3383 3 1 3457 XNOR3X2 $T=1123980 866320 0 0 $X=1123978 $Y=865918
X913 3570 3453 3457 3 1 3844 XNOR3X2 $T=1149060 856240 1 0 $X=1149058 $Y=850800
X914 3687 3645 3507 3 1 3661 XNOR3X2 $T=1183380 886480 1 180 $X=1171500 $Y=886078
X915 3867 3593 3845 3 1 4047 XNOR3X2 $T=1206480 926800 1 0 $X=1206478 $Y=921360
X916 3448 3871 3848 3 1 4028 XNOR3X2 $T=1219680 755440 0 0 $X=1219678 $Y=755038
X917 4091 4047 4170 3 1 4173 XNOR3X2 $T=1242120 926800 0 0 $X=1242118 $Y=926398
X918 3936 4219 4110 3 1 4278 XNOR3X2 $T=1265880 946960 0 0 $X=1265878 $Y=946558
X919 4414 4359 4381 3 1 4496 XNOR3X2 $T=1307460 765520 0 0 $X=1307458 $Y=765118
X920 2504 1 2505 2478 2366 2397 3 AOI22XL $T=916080 946960 1 180 $X=912780 $Y=946558
X921 2799 1 2780 2864 2865 2736 3 AOI22XL $T=991320 926800 0 0 $X=991318 $Y=926398
X922 188 1 6066 6050 183 6002 3 AOI22XL $T=1644060 896560 0 180 $X=1640760 $Y=891120
X923 185 1 6066 6050 188 6003 3 AOI22XL $T=1646040 896560 1 180 $X=1642740 $Y=896158
X924 193 1 6046 189 188 6059 3 AOI22XL $T=1646040 957040 0 180 $X=1642740 $Y=951600
X925 193 1 6118 189 183 6067 3 AOI22XL $T=1653960 957040 0 180 $X=1650660 $Y=951600
X926 193 1 6185 189 184 6126 3 AOI22XL $T=1659240 936880 0 180 $X=1655940 $Y=931440
X927 194 1 6066 6050 190 6159 3 AOI22XL $T=1661220 896560 1 0 $X=1661218 $Y=891120
X928 190 1 6066 6050 184 6027 3 AOI22XL $T=1664520 886480 1 180 $X=1661220 $Y=886078
X929 198 1 6066 6050 185 6142 3 AOI22XL $T=1672440 896560 0 180 $X=1669140 $Y=891120
X930 184 1 6066 6050 199 6204 3 AOI22XL $T=1671780 886480 0 0 $X=1671778 $Y=886078
X931 193 1 6160 189 190 6207 3 AOI22XL $T=1671780 957040 1 0 $X=1671778 $Y=951600
X932 193 1 6208 189 199 6226 3 AOI22XL $T=1674420 936880 0 0 $X=1674418 $Y=936478
X933 199 1 6066 6050 202 6249 3 AOI22XL $T=1684320 896560 1 0 $X=1684318 $Y=891120
X934 202 1 6066 6050 203 6373 3 AOI22XL $T=1709400 896560 0 180 $X=1706100 $Y=891120
X935 193 1 6316 189 202 6422 3 AOI22XL $T=1709400 936880 1 0 $X=1709398 $Y=931440
X936 193 1 6368 189 203 6405 3 AOI22XL $T=1710720 946960 0 0 $X=1710718 $Y=946558
X937 193 1 6369 189 210 6420 3 AOI22XL $T=1712040 977200 1 0 $X=1712038 $Y=971760
X938 203 1 6066 6050 210 6429 3 AOI22XL $T=1717320 896560 0 0 $X=1717318 $Y=896158
X939 210 1 6066 6050 212 6428 3 AOI22XL $T=1718640 906640 0 0 $X=1718638 $Y=906238
X940 205 1 199 203 202 201 3 NOR4BX1 $T=1685640 967120 1 180 $X=1681680 $Y=966718
X941 6406 213 3 1 BUFX4 $T=1714680 836080 0 0 $X=1714678 $Y=835678
X942 7622 7649 3 1 7616 NAND2BX4 $T=1976700 957040 1 0 $X=1976698 $Y=951600
X943 8112 8072 3 1 7941 NAND2BX4 $T=2073720 826000 1 180 $X=2068440 $Y=825598
X944 203 207 210 1 3 350 OR3XL $T=1695540 977200 1 180 $X=1692240 $Y=976798
X945 7901 3 7834 1 7810 7875 NAND3XL $T=2024880 957040 1 180 $X=2022240 $Y=956638
X946 7880 3 7939 1 7971 7976 NAND3XL $T=2042040 826000 0 0 $X=2042038 $Y=825598
X947 7971 3 7941 1 8092 8056 NAND3XL $T=2068440 805840 0 0 $X=2068438 $Y=805438
X948 4174 4077 3155 3 4186 1 OAI2BB1XL $T=1256640 775600 0 0 $X=1256638 $Y=775198
X949 7131 7108 224 1 3 7190 NAND3BX2 $T=1877040 957040 1 0 $X=1877038 $Y=951600
X950 3623 3379 3 3619 1 3614 3617 OAI211XL $T=1164900 775600 1 180 $X=1160940 $Y=775198
X951 180 179 183 6035 173 1 3 188 SDFFRHQX1 $T=1633500 926800 1 0 $X=1633498 $Y=921360
X952 180 179 188 6091 173 1 3 184 SDFFRHQX1 $T=1653960 916720 0 180 $X=1637460 $Y=911280
X953 180 179 194 6161 173 1 3 190 SDFFRHQX1 $T=1668480 967120 1 180 $X=1651980 $Y=966718
X954 180 179 184 6194 173 1 3 199 SDFFRHQX1 $T=1667160 916720 1 0 $X=1667158 $Y=911280
X955 180 179 203 6423 173 1 3 210 SDFFRHQX1 $T=1713360 967120 1 0 $X=1713358 $Y=961680
X956 180 179 202 6462 173 1 3 203 SDFFRHQX1 $T=1730520 936880 1 180 $X=1714020 $Y=936478
X957 180 179 214 6426 173 1 3 202 SDFFRHQX1 $T=1714680 916720 1 0 $X=1714678 $Y=911280
X958 3875 3 3842 3763 3719 3843 1 NAND4X1 $T=1203840 826000 1 180 $X=1200540 $Y=825598
X959 7877 3 7977 247 7969 7946 1 NAND4X1 $T=2045340 926800 0 180 $X=2042040 $Y=921360
X960 8051 3 8049 7939 1 8072 NAND3X4 $T=2062500 856240 0 180 $X=2055900 $Y=850800
X961 4053 3 4107 4130 1 4046 NAND3BX1 $T=1250040 896560 0 180 $X=1246740 $Y=891120
X962 3843 3998 3 4010 3843 3747 1 3841 OAI221X2 $T=1226940 826000 1 0 $X=1226938 $Y=820560
X963 82 3462 3483 3482 3 1 MXI2X2 $T=1137180 946960 1 0 $X=1137178 $Y=941520
X964 4213 4188 3 4196 4194 4381 1 AOI2BB2X2 $T=1263240 765520 0 0 $X=1263238 $Y=765118
X965 3844 3801 3763 1 3866 3725 3850 3 AOI32X2 $T=1202520 846160 1 0 $X=1202518 $Y=840720
X966 199 202 203 204 3 1 351 AND4X2 $T=1684320 977200 0 0 $X=1684318 $Y=976798
X967 7896 7855 7809 7853 7405 1 3 OAI31X4 $T=2022240 866320 1 180 $X=2016300 $Y=865918
X968 7941 7927 7897 7926 7232 1 3 OAI31X4 $T=2036760 815920 1 180 $X=2030820 $Y=815518
X969 8057 7948 1 8073 8050 3 7833 NAND4X2 $T=2063820 846160 0 180 $X=2057880 $Y=840720
X970 8089 8141 8138 8004 8146 1 7794 3 OAI32X4 $T=2079000 815920 1 0 $X=2078998 $Y=810480
.ENDS
***************************************
.SUBCKT OAI222X2 B1 B0 VSS A0 A1 C0 C1 Y VDD
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4BXL AN VDD D C B Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDFX1 B A CI CO VSS VDD S
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_63 2 4 26 27 28 29 31 34 35 37 38 39 41 42 43 44 45 46 47 48
+ 49 50 51 52 53 54 55 56 57 58 59 60 61 63 65 67 68 69 71 72
+ 73 75 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94
+ 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114
+ 115 116 117 118 119 120 122 123 125 126 127 129 131 132 133 134 136 137 138 140
+ 141 142 143 144 145 147 148 149 151 152 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205
+ 206 207 211 212 213 214 215 217 218 219 220 221 222 223 224 225 226 227 228 229
+ 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 250
+ 251 252 253 254 255 256 257 258 259 260 261 262 263 264 265 266 267 268 269 270
+ 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286 287 288 289 290
+ 291 292 293 294 295 296 297 298 299 300 301 302 303 304 305 306 307 308 309 310
+ 311 312 313 314 315 316 317 318 319 320 322 323 324 325 326 327 329 330 332 333
+ 334 335 337 338 339 340 341 342 343 345 347 348 350 352 353 354 355 356 358 359
+ 361 362 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381
+ 382 383 384 385 386 387 388 389 390 391 392 394 395 396 398 399 400 401 402 403
+ 404 405 406 407 408 409 410 411 412 413 414 416 417 418 419 420 421 422 423 424
+ 427 428 429 431 433 438 440 442 444 445 446 451 452 453 454 455 456 1267 1268
** N=23502 EP=379 IP=6647 FDC=0
X0 1591 4 1578 2 1601 NAND2X1 $T=772860 1108240 1 180 $X=770880 $Y=1107838
X1 37 4 1698 2 1713 NAND2X1 $T=805200 1108240 0 0 $X=805198 $Y=1107838
X2 1577 4 1776 2 1774 NAND2X1 $T=834900 1027600 0 0 $X=834898 $Y=1027198
X3 1715 4 1777 2 1795 NAND2X1 $T=836220 1057840 1 0 $X=836218 $Y=1052400
X4 1685 4 1778 2 1805 NAND2X1 $T=844140 1078000 1 180 $X=842160 $Y=1077598
X5 57 4 56 2 2019 NAND2X1 $T=927300 1108240 0 180 $X=925320 $Y=1102800
X6 59 4 58 2 2037 NAND2X1 $T=938520 1098160 0 0 $X=938518 $Y=1097758
X7 61 4 60 2 2046 NAND2X1 $T=941820 1128400 0 180 $X=939840 $Y=1122960
X8 2175 4 2176 2 2160 NAND2X1 $T=958980 1078000 0 180 $X=957000 $Y=1072560
X9 2209 4 2161 2 2162 NAND2X1 $T=969540 1017520 0 180 $X=967560 $Y=1012080
X10 2222 4 69 2 2114 NAND2X1 $T=974160 1138480 1 0 $X=974158 $Y=1133040
X11 2206 4 2209 2 2233 NAND2X1 $T=976800 987280 0 0 $X=976798 $Y=986878
X12 2283 4 2267 2 2282 NAND2X1 $T=991320 1027600 0 180 $X=989340 $Y=1022160
X13 2267 4 2268 2 2163 NAND2X1 $T=991320 1037680 0 180 $X=989340 $Y=1032240
X14 2251 4 2287 2 2174 NAND2X1 $T=994620 997360 0 0 $X=994618 $Y=996958
X15 72 4 2286 2 2206 NAND2X1 $T=995940 987280 1 0 $X=995938 $Y=981840
X16 2278 4 2197 2 2321 NAND2X1 $T=998580 1088080 1 0 $X=998578 $Y=1082640
X17 2288 4 2339 2 2341 NAND2X1 $T=1006500 1088080 0 0 $X=1006498 $Y=1087678
X18 2385 4 2360 2 2322 NAND2X1 $T=1015740 1037680 1 180 $X=1013760 $Y=1037278
X19 2358 4 2359 2 2283 NAND2X1 $T=1019700 1017520 0 0 $X=1019698 $Y=1017118
X20 2477 4 2381 2 2281 NAND2X1 $T=1021680 1088080 0 180 $X=1019700 $Y=1082640
X21 2389 4 2388 2 2335 NAND2X1 $T=1025640 1067920 0 180 $X=1023660 $Y=1062480
X22 2416 4 2414 2 2386 NAND2X1 $T=1034880 1138480 0 180 $X=1032900 $Y=1133040
X23 85 4 2448 2 82 NAND2X1 $T=1048740 1138480 0 180 $X=1046760 $Y=1133040
X24 2561 4 2591 2 2551 NAND2X1 $T=1094280 1118320 0 0 $X=1094278 $Y=1117918
X25 145 4 2841 2 151 NAND2X1 $T=1228920 1118320 0 0 $X=1228918 $Y=1117918
X26 2988 4 151 2 3046 NAND2X1 $T=1242120 1118320 0 0 $X=1242118 $Y=1117918
X27 3104 4 3110 2 3141 NAND2X1 $T=1247400 1037680 1 0 $X=1247398 $Y=1032240
X28 3199 4 3152 2 3209 NAND2X1 $T=1275780 1088080 0 0 $X=1275778 $Y=1087678
X29 179 4 182 2 184 NAND2X1 $T=1383360 987280 0 0 $X=1383358 $Y=986878
X30 3557 4 3595 2 3621 NAND2X1 $T=1427580 1118320 0 0 $X=1427578 $Y=1117918
X31 194 4 3596 2 3653 NAND2X1 $T=1435500 1128400 0 0 $X=1435498 $Y=1127998
X32 3582 4 3606 2 3759 NAND2X1 $T=1461900 1088080 0 0 $X=1461898 $Y=1087678
X33 3604 4 3713 2 3775 NAND2X1 $T=1465200 1067920 1 0 $X=1465198 $Y=1062480
X34 3635 4 3724 2 3786 NAND2X1 $T=1470480 1017520 1 0 $X=1470478 $Y=1012080
X35 3759 4 3756 2 3792 NAND2X1 $T=1478400 1088080 0 0 $X=1478398 $Y=1087678
X36 3788 4 3793 2 3823 NAND2X1 $T=1485000 1118320 0 0 $X=1484998 $Y=1117918
X37 3775 4 3714 2 3808 NAND2X1 $T=1490280 1067920 1 0 $X=1490278 $Y=1062480
X38 3463 4 3908 2 3957 NAND2X1 $T=1521960 1057840 1 180 $X=1519980 $Y=1057438
X39 3451 4 3909 2 3971 NAND2X1 $T=1525920 1088080 1 0 $X=1525918 $Y=1082640
X40 3942 4 3920 2 4051 NAND2X1 $T=1551660 1057840 1 180 $X=1549680 $Y=1057438
X41 3317 4 4038 2 4053 NAND2X1 $T=1560900 1007440 0 0 $X=1560898 $Y=1007038
X42 4104 4 1875 2 4137 NAND2X1 $T=1582020 1047760 0 0 $X=1582018 $Y=1047358
X43 223 4 219 2 218 NAND2X1 $T=1622280 1057840 0 0 $X=1622278 $Y=1057438
X44 4384 4 4326 2 4381 NAND2X1 $T=1641420 1088080 0 180 $X=1639440 $Y=1082640
X45 4381 4 4388 2 4411 NAND2X1 $T=1663860 1088080 1 0 $X=1663858 $Y=1082640
X46 4342 4 4482 2 4481 NAND2X1 $T=1688940 1108240 0 0 $X=1688938 $Y=1107838
X47 4574 4 4573 2 4589 NAND2X1 $T=1712700 1098160 1 180 $X=1710720 $Y=1097758
X48 261 4 259 2 4572 NAND2X1 $T=1714680 1128400 1 180 $X=1712700 $Y=1127998
X49 262 4 259 2 4604 NAND2X1 $T=1722600 1128400 1 180 $X=1720620 $Y=1127998
X50 4787 4 3929 2 4742 NAND2X1 $T=1760880 1108240 1 180 $X=1758900 $Y=1107838
X51 4782 4 4267 2 4756 NAND2X1 $T=1764180 1017520 1 180 $X=1762200 $Y=1017118
X52 4806 4 4088 2 4770 NAND2X1 $T=1772100 1098160 1 180 $X=1770120 $Y=1097758
X53 4783 4 4831 2 4804 NAND2X1 $T=1778040 1057840 0 0 $X=1778038 $Y=1057438
X54 4818 4 4269 2 266 NAND2X1 $T=1783320 997360 0 180 $X=1781340 $Y=991920
X55 4788 4 4808 2 4853 NAND2X1 $T=1793220 1098160 0 0 $X=1793218 $Y=1097758
X56 4831 4 4801 2 4864 NAND2X1 $T=1793880 1007440 0 0 $X=1793878 $Y=1007038
X57 273 4 4922 2 4923 NAND2X1 $T=1809720 1037680 1 0 $X=1809718 $Y=1032240
X58 276 4 4964 2 4982 NAND2X1 $T=1828860 1057840 0 0 $X=1828858 $Y=1057438
X59 278 4 4976 2 4980 NAND2X1 $T=1831500 1047760 0 0 $X=1831498 $Y=1047358
X60 5007 4 5006 2 289 NAND2X1 $T=1845360 1078000 0 180 $X=1843380 $Y=1072560
X61 292 4 293 2 5086 NAND2X1 $T=1867140 1118320 1 0 $X=1867138 $Y=1112880
X62 294 4 5118 2 5083 NAND2X1 $T=1872420 1047760 1 0 $X=1872418 $Y=1042320
X63 5131 4 5138 2 297 NAND2X1 $T=1877700 987280 0 0 $X=1877698 $Y=986878
X64 303 4 5172 2 5182 NAND2X1 $T=1888260 1037680 1 0 $X=1888258 $Y=1032240
X65 5267 4 5051 2 305 NAND2X1 $T=1892220 1057840 1 180 $X=1890240 $Y=1057438
X66 308 4 5244 2 5245 NAND2X1 $T=1906080 1047760 1 0 $X=1906078 $Y=1042320
X67 314 4 5286 2 5354 NAND2X1 $T=1919280 1027600 1 0 $X=1919278 $Y=1022160
X68 319 4 5328 2 5323 NAND2X1 $T=1929840 1037680 1 0 $X=1929838 $Y=1032240
X69 323 4 322 2 5303 NAND2X1 $T=1943040 1108240 0 180 $X=1941060 $Y=1102800
X70 326 4 325 2 5424 NAND2X1 $T=1956240 1118320 0 0 $X=1956238 $Y=1117918
X71 334 4 335 2 5483 NAND2X1 $T=2003100 1138480 1 0 $X=2003098 $Y=1133040
X72 5596 4 5564 2 5583 NAND2X1 $T=2020920 1088080 1 180 $X=2018940 $Y=1087678
X73 5592 4 5594 2 5623 NAND2X1 $T=2038740 1067920 0 0 $X=2038738 $Y=1067518
X74 340 4 343 2 5641 NAND2X1 $T=2046660 1138480 1 0 $X=2046658 $Y=1133040
X75 5767 4 5714 2 5628 NAND2X1 $T=2059200 1098160 0 0 $X=2059198 $Y=1097758
X76 5728 4 5758 2 5772 NAND2X1 $T=2066460 987280 0 0 $X=2066458 $Y=986878
X77 5771 4 5773 2 5679 NAND2X1 $T=2075040 1057840 1 0 $X=2075038 $Y=1052400
X78 5802 4 5801 2 5726 NAND2X1 $T=2084940 1007440 1 180 $X=2082960 $Y=1007038
X79 5832 4 5830 2 5742 NAND2X1 $T=2096160 1027600 1 180 $X=2094180 $Y=1027198
X80 5798 4 5831 2 342 NAND2X1 $T=2094840 997360 0 0 $X=2094838 $Y=996958
X81 5893 4 5891 2 5798 NAND2X1 $T=2107380 997360 0 0 $X=2107378 $Y=996958
X82 6185 4 6149 2 395 NAND2X1 $T=2203740 997360 1 0 $X=2203738 $Y=991920
X83 6230 4 383 2 6350 NAND2X1 $T=2264460 1057840 0 0 $X=2264458 $Y=1057438
X84 6410 4 6509 2 6510 NAND2X1 $T=2325180 1108240 0 0 $X=2325178 $Y=1107838
X85 6363 4 6452 2 6563 NAND2X1 $T=2343000 1128400 1 0 $X=2342998 $Y=1122960
X86 6525 4 6486 2 6593 NAND2X1 $T=2356200 1098160 1 0 $X=2356198 $Y=1092720
X87 6640 4 422 2 6702 NAND2X1 $T=2387220 1118320 0 0 $X=2387218 $Y=1117918
X88 6687 4 6730 2 6739 NAND2X1 $T=2403060 1098160 1 0 $X=2403058 $Y=1092720
X89 7015 4 7002 2 7001 NAND2X1 $T=2504040 1118320 0 180 $X=2502060 $Y=1112880
X90 446 4 445 2 7015 NAND2X1 $T=2511300 1128400 1 180 $X=2509320 $Y=1127998
X91 7149 4 451 2 7090 NAND2X1 $T=2543640 1118320 0 180 $X=2541660 $Y=1112880
X92 37 2 4 1698 1714 NOR2X4 $T=815100 1108240 1 180 $X=810480 $Y=1107838
X93 3704 2 4 3638 3807 NOR2X4 $T=1485000 1037680 1 0 $X=1484998 $Y=1032240
X94 3366 2 4 3986 4008 NOR2X4 $T=1549680 1027600 1 180 $X=1545060 $Y=1027198
X95 211 2 4 1877 4106 NOR2X4 $T=1577400 1118320 1 180 $X=1572780 $Y=1117918
X96 4360 2 4 4339 4382 NOR2X4 $T=1654620 1108240 1 180 $X=1650000 $Y=1107838
X97 4419 2 4 4382 4426 NOR2X4 $T=1671120 1108240 0 0 $X=1671118 $Y=1107838
X98 4771 2 4 4087 4773 NOR2X4 $T=1772100 1057840 0 180 $X=1767480 $Y=1052400
X99 2038 4 2046 53 2 NAND2BX1 $T=918720 1128400 1 180 $X=916080 $Y=1127998
X100 1983 4 2019 1976 2 NAND2BX1 $T=922680 1108240 0 180 $X=920040 $Y=1102800
X101 2062 4 2037 1958 2 NAND2BX1 $T=927960 1098160 1 180 $X=925320 $Y=1097758
X102 2411 4 2386 2365 2 NAND2BX1 $T=1024320 1138480 0 180 $X=1021680 $Y=1133040
X103 111 4 2674 122 2 NAND2BX1 $T=1127940 987280 1 0 $X=1127938 $Y=981840
X104 3167 4 3143 3176 2 NAND2BX1 $T=1265880 1007440 1 0 $X=1265878 $Y=1002000
X105 3702 4 3653 195 2 NAND2BX1 $T=1450680 1128400 0 0 $X=1450678 $Y=1127998
X106 3725 4 3621 3747 2 NAND2BX1 $T=1469160 1128400 1 0 $X=1469158 $Y=1122960
X107 3729 4 3786 3803 2 NAND2BX1 $T=1482360 1027600 1 0 $X=1482358 $Y=1022160
X108 3807 4 3773 3867 2 NAND2BX1 $T=1503480 1037680 1 0 $X=1503478 $Y=1032240
X109 4008 4 4060 4223 2 NAND2BX1 $T=1595880 1027600 0 0 $X=1595878 $Y=1027198
X110 5578 4 5564 5563 2 NAND2BX1 $T=2015640 1088080 1 180 $X=2013000 $Y=1087678
X111 5681 4 5679 5667 2 NAND2BX1 $T=2047980 1027600 0 180 $X=2045340 $Y=1022160
X112 5727 4 5726 5713 2 NAND2BX1 $T=2057880 997360 1 180 $X=2055240 $Y=996958
X113 5729 4 5742 5626 2 NAND2BX1 $T=2063820 1027600 1 0 $X=2063818 $Y=1022160
X114 6536 4 6510 421 2 NAND2BX1 $T=2346960 1118320 0 0 $X=2346958 $Y=1117918
X115 6775 4 6776 6834 2 NAND2BX1 $T=2439360 1118320 0 0 $X=2439358 $Y=1117918
X116 1775 1850 4 1805 2 1876 OAI21X1 $T=852060 1067920 0 0 $X=852058 $Y=1067518
X117 2038 54 4 2046 2 2007 OAI21X1 $T=916080 1128400 1 0 $X=916078 $Y=1122960
X118 2325 67 4 2320 2 2280 OAI21X1 $T=1002540 1067920 0 180 $X=999240 $Y=1062480
X119 3702 197 4 3653 2 3743 OAI21X1 $T=1457280 1128400 0 0 $X=1457278 $Y=1127998
X120 3653 3725 4 3621 2 3733 OAI21X1 $T=1463880 1128400 1 0 $X=1463878 $Y=1122960
X121 3773 3729 4 3786 2 3789 OAI21X1 $T=1488300 1017520 1 180 $X=1485000 $Y=1017118
X122 4864 4817 4 4790 2 4863 OAI21X1 $T=1800480 1007440 0 180 $X=1797180 $Y=1002000
X123 5607 5608 4 5623 2 5639 OAI21X1 $T=2031480 1067920 1 0 $X=2031478 $Y=1062480
X124 6624 424 4 6564 2 423 OAI21X1 $T=2373360 1138480 0 180 $X=2370060 $Y=1133040
X125 6704 424 4 6677 2 6691 OAI21X1 $T=2399100 1128400 1 180 $X=2395800 $Y=1127998
X126 1805 4 1790 1795 2 1804 OAI21XL $T=844800 1067920 0 180 $X=842160 $Y=1062480
X127 2062 4 2019 2037 2 2034 OAI21XL $T=917400 1098160 1 180 $X=914760 $Y=1097758
X128 2163 4 2187 2189 2 2190 OAI21XL $T=958980 1037680 0 0 $X=958978 $Y=1037278
X129 67 4 2191 2192 2 2158 OAI21XL $T=962940 1067920 0 180 $X=960300 $Y=1062480
X130 2162 4 2189 2195 2 2193 OAI21XL $T=961620 1027600 1 0 $X=961618 $Y=1022160
X131 2205 4 2160 2194 2 2173 OAI21XL $T=964260 1088080 0 180 $X=961620 $Y=1082640
X132 2187 4 2220 2218 2 2226 OAI21XL $T=972180 1037680 0 0 $X=972178 $Y=1037278
X133 2219 4 67 2225 2 2231 OAI21XL $T=973500 1067920 1 0 $X=973498 $Y=1062480
X134 2114 4 67 2205 2 2250 OAI21XL $T=973500 1108240 1 0 $X=973498 $Y=1102800
X135 2281 4 2330 2335 2 2234 OAI21XL $T=1003200 1078000 1 0 $X=1003198 $Y=1072560
X136 82 4 2411 2386 2 2295 OAI21XL $T=1040160 1138480 0 180 $X=1037520 $Y=1133040
X137 109 4 107 105 2 113 OAI21XL $T=1129260 1037680 0 180 $X=1126620 $Y=1032240
X138 102 4 94 91 2 2674 OAI21XL $T=1130580 1017520 0 180 $X=1127940 $Y=1012080
X139 115 4 96 102 2 2710 OAI21XL $T=1137180 1067920 1 0 $X=1137178 $Y=1062480
X140 120 4 119 103 2 2850 OAI21XL $T=1176120 1098160 0 0 $X=1176118 $Y=1097758
X141 2786 4 2795 2823 2 2835 OAI21XL $T=1176780 997360 1 0 $X=1176778 $Y=991920
X142 108 4 110 104 2 2839 OAI21XL $T=1177440 1067920 1 0 $X=1177438 $Y=1062480
X143 119 4 107 2836 2 2885 OAI21XL $T=1180080 1017520 0 0 $X=1180078 $Y=1017118
X144 88 4 91 104 2 2836 OAI21XL $T=1180080 1027600 0 0 $X=1180078 $Y=1027198
X145 2849 4 2841 2839 2 132 OAI21XL $T=1186680 1067920 0 180 $X=1184040 $Y=1062480
X146 88 4 136 2850 2 133 OAI21XL $T=1190640 1098160 1 180 $X=1188000 $Y=1097758
X147 2849 4 100 137 2 2873 OAI21XL $T=1193280 1067920 1 0 $X=1193278 $Y=1062480
X148 110 4 96 2873 2 2989 OAI21XL $T=1194600 1047760 0 0 $X=1194598 $Y=1047358
X149 141 4 2849 102 2 2947 OAI21XL $T=1209120 1088080 0 180 $X=1206480 $Y=1082640
X150 145 4 120 2978 2 2972 OAI21XL $T=1219680 1108240 1 180 $X=1217040 $Y=1107838
X151 145 4 2841 115 2 2988 OAI21XL $T=1219680 1118320 1 180 $X=1217040 $Y=1117918
X152 136 4 129 95 2 2978 OAI21XL $T=1219680 1128400 0 180 $X=1217040 $Y=1122960
X153 147 4 2799 2989 2 3027 OAI21XL $T=1229580 1037680 0 180 $X=1226940 $Y=1032240
X154 149 4 3049 3051 2 3069 OAI21XL $T=1232220 1067920 1 0 $X=1232218 $Y=1062480
X155 3046 4 148 88 2 3045 OAI21XL $T=1234860 1078000 1 180 $X=1232220 $Y=1077598
X156 3047 4 3068 3027 2 3154 OAI21XL $T=1237500 1027600 0 0 $X=1237498 $Y=1027198
X157 152 4 3090 2971 2 3142 OAI21XL $T=1242780 1088080 1 0 $X=1242778 $Y=1082640
X158 3118 4 3105 3140 2 3199 OAI21XL $T=1255980 1108240 0 0 $X=1255978 $Y=1107838
X159 3177 4 3144 3141 2 3169 OAI21XL $T=1267860 1037680 0 180 $X=1265220 $Y=1032240
X160 3245 4 3195 3177 2 3242 OAI21XL $T=1291620 1047760 1 180 $X=1288980 $Y=1047358
X161 5260 4 5235 5249 2 5300 OAI21XL $T=1922580 1088080 1 0 $X=1922578 $Y=1082640
X162 5583 4 5597 5608 2 5613 OAI21XL $T=2024880 1088080 1 0 $X=2024878 $Y=1082640
X163 5643 4 5597 5628 2 5580 OAI21XL $T=2039400 1108240 0 180 $X=2036760 $Y=1102800
X164 5727 4 5744 5726 2 5684 OAI21XL $T=2067120 1007440 1 180 $X=2064480 $Y=1007038
X165 5793 4 5726 5798 2 5788 OAI21XL $T=2080980 997360 0 0 $X=2080978 $Y=996958
X166 6563 4 6536 6510 2 6621 OAI21XL $T=2346960 1108240 0 0 $X=2346958 $Y=1107838
X167 6593 4 6610 6609 2 6611 OAI21XL $T=2364780 1098160 1 0 $X=2364778 $Y=1092720
X168 6636 4 6677 6674 2 6675 OAI21XL $T=2392500 1108240 1 180 $X=2389860 $Y=1107838
X169 6739 4 424 6676 2 6742 OAI21XL $T=2408340 1098160 1 0 $X=2408338 $Y=1092720
X170 6741 4 424 6688 2 6740 OAI21XL $T=2408340 1098160 0 0 $X=2408338 $Y=1097758
X171 6702 4 424 6703 2 6774 OAI21XL $T=2414280 1118320 0 0 $X=2414278 $Y=1117918
X172 6775 4 6703 6776 2 431 OAI21XL $T=2423520 1128400 1 0 $X=2423518 $Y=1122960
X173 1821 1850 1877 4 2 XOR2X4 $T=847440 1098160 1 0 $X=847438 $Y=1092720
X174 1756 1861 1874 4 2 XOR2X4 $T=848760 1118320 0 0 $X=848758 $Y=1117918
X175 1849 1876 1901 4 2 XOR2X4 $T=862620 1067920 0 0 $X=862618 $Y=1067518
X176 4009 4037 4088 4 2 XOR2X4 $T=1548360 1098160 1 0 $X=1548358 $Y=1092720
X177 4169 4198 4269 4 2 XOR2X4 $T=1593240 1007440 0 0 $X=1593238 $Y=1007038
X178 4220 4235 4265 4 2 XOR2X4 $T=1602480 1047760 0 0 $X=1602478 $Y=1047358
X179 4234 217 4418 4 2 XOR2X4 $T=1614360 1118320 0 0 $X=1614358 $Y=1117918
X180 4151 4249 4339 4 2 XOR2X4 $T=1617660 1108240 0 0 $X=1617658 $Y=1107838
X181 5626 5612 5492 4 2 XOR2X4 $T=2036100 1027600 0 180 $X=2024880 $Y=1022160
X182 442 6944 4594 4 2 XOR2X4 $T=2493480 1108240 0 180 $X=2482260 $Y=1102800
X183 1639 4 2 1605 INVX1 $T=786060 1118320 1 180 $X=784740 $Y=1117918
X184 1714 4 2 1729 INVX1 $T=814440 1118320 1 180 $X=813120 $Y=1117918
X185 1804 4 2 1803 INVX1 $T=842820 1057840 0 180 $X=841500 $Y=1052400
X186 51 4 2 43 INVX1 $T=908820 987280 0 180 $X=907500 $Y=981840
X187 1983 4 2 2032 INVX1 $T=914100 1108240 1 180 $X=912780 $Y=1107838
X188 2174 4 2 2217 INVX1 $T=959640 1007440 1 0 $X=959638 $Y=1002000
X189 2206 4 2 2207 INVX1 $T=967560 997360 1 0 $X=967558 $Y=991920
X190 2234 4 2 2187 INVX1 $T=979440 1037680 1 180 $X=978120 $Y=1037278
X191 2249 4 2 2189 INVX1 $T=982080 1027600 0 180 $X=980760 $Y=1022160
X192 2322 4 2 2294 INVX1 $T=999240 1027600 1 180 $X=997920 $Y=1027198
X193 92 4 2 94 INVX1 $T=1078440 987280 1 0 $X=1078438 $Y=981840
X194 110 4 2 2558 INVX1 $T=1121340 1047760 0 180 $X=1120020 $Y=1042320
X195 89 4 2 109 INVX1 $T=1138500 997360 1 180 $X=1137180 $Y=996958
X196 2726 4 2 2714 INVX1 $T=1147080 1027600 0 180 $X=1145760 $Y=1022160
X197 2797 4 2 2784 INVX1 $T=1167540 1027600 0 180 $X=1166220 $Y=1022160
X198 110 4 2 2849 INVX1 $T=1178100 1078000 0 180 $X=1176780 $Y=1072560
X199 108 4 2 2841 INVX1 $T=1186020 1118320 1 180 $X=1184700 $Y=1117918
X200 2885 4 2 3017 INVX1 $T=1224960 1007440 0 0 $X=1224958 $Y=1007038
X201 2799 4 2 3047 INVX1 $T=1231560 1027600 0 0 $X=1231558 $Y=1027198
X202 147 4 2 3068 INVX1 $T=1234200 1037680 0 0 $X=1234198 $Y=1037278
X203 3091 4 2 3143 INVX1 $T=1243440 1007440 1 0 $X=1243438 $Y=1002000
X204 3154 4 2 3192 INVX1 $T=1260600 1017520 0 0 $X=1260598 $Y=1017118
X205 3169 4 2 3167 INVX1 $T=1268520 1027600 0 180 $X=1267200 $Y=1022160
X206 3144 4 2 3211 INVX1 $T=1273800 1037680 1 0 $X=1273798 $Y=1032240
X207 3305 4 2 3451 INVX1 $T=1320660 1088080 0 0 $X=1320658 $Y=1087678
X208 3775 4 2 3770 INVX1 $T=1481700 1067920 0 180 $X=1480380 $Y=1062480
X209 3295 4 2 3788 INVX1 $T=1483020 1128400 0 0 $X=1483018 $Y=1127998
X210 3890 4 2 206 INVX1 $T=1511400 1128400 0 0 $X=1511398 $Y=1127998
X211 3957 4 2 3989 INVX1 $T=1535160 1057840 0 0 $X=1535158 $Y=1057438
X212 4172 4 2 4104 INVX1 $T=1593900 1057840 0 180 $X=1592580 $Y=1052400
X213 4103 4 2 4194 INVX1 $T=1595220 1078000 0 0 $X=1595218 $Y=1077598
X214 4161 4 2 4236 INVX1 $T=1605780 1098160 0 0 $X=1605778 $Y=1097758
X215 4405 4 2 4410 INVX1 $T=1663200 997360 0 0 $X=1663198 $Y=996958
X216 4406 4 2 4442 INVX1 $T=1663200 1037680 1 0 $X=1663198 $Y=1032240
X217 4404 4 2 4446 INVX1 $T=1665840 1098160 1 0 $X=1665838 $Y=1092720
X218 4434 4 2 239 INVX1 $T=1679040 1007440 1 0 $X=1679038 $Y=1002000
X219 4382 4 2 4482 INVX1 $T=1681680 1108240 0 0 $X=1681678 $Y=1107838
X220 245 4 2 4420 INVX1 $T=1685640 1007440 1 180 $X=1684320 $Y=1007038
X221 255 4 2 256 INVX1 $T=1698840 1007440 1 0 $X=1698838 $Y=1002000
X222 4564 4 2 4600 INVX1 $T=1708080 1027600 0 0 $X=1708078 $Y=1027198
X223 4575 4 2 4592 INVX1 $T=1713360 1007440 0 0 $X=1713358 $Y=1007038
X224 4577 4 2 4606 INVX1 $T=1723260 987280 0 0 $X=1723258 $Y=986878
X225 4756 4 2 4789 INVX1 $T=1768140 1017520 1 0 $X=1768138 $Y=1012080
X226 4770 4 2 4772 INVX1 $T=1768140 1088080 0 0 $X=1768138 $Y=1087678
X227 4742 4 2 4821 INVX1 $T=1781340 1128400 1 0 $X=1781338 $Y=1122960
X228 4773 4 2 4831 INVX1 $T=1788600 1047760 0 0 $X=1788598 $Y=1047358
X229 4974 4 2 4978 INVX1 $T=1830840 1128400 1 0 $X=1830838 $Y=1122960
X230 4994 4 2 4981 INVX1 $T=1840080 1088080 1 180 $X=1838760 $Y=1087678
X231 5064 4 2 5066 INVX1 $T=1857900 1067920 1 0 $X=1857898 $Y=1062480
X232 5086 4 2 5099 INVX1 $T=1865160 1118320 0 180 $X=1863840 $Y=1112880
X233 5141 4 2 5082 INVX1 $T=1880340 1047760 0 180 $X=1879020 $Y=1042320
X234 298 4 2 5133 INVX1 $T=1880340 1128400 1 0 $X=1880338 $Y=1122960
X235 302 4 2 5084 INVX1 $T=1883640 1098160 1 180 $X=1882320 $Y=1097758
X236 5195 4 2 5203 INVX1 $T=1896180 1057840 1 0 $X=1896178 $Y=1052400
X237 5193 4 2 5235 INVX1 $T=1896180 1098160 1 0 $X=1896178 $Y=1092720
X238 5289 4 2 327 INVX1 $T=1930500 1138480 1 0 $X=1930498 $Y=1133040
X239 5327 4 2 5295 INVX1 $T=1932480 1057840 0 0 $X=1932478 $Y=1057438
X240 5336 4 2 5367 INVX1 $T=1941720 1057840 1 0 $X=1941718 $Y=1052400
X241 312 4 2 329 INVX1 $T=1950960 1138480 1 0 $X=1950958 $Y=1133040
X242 5399 4 2 330 INVX1 $T=1957560 1138480 0 180 $X=1956240 $Y=1133040
X243 5424 4 2 5427 INVX1 $T=1969440 1118320 0 0 $X=1969438 $Y=1117918
X244 5310 4 2 5425 INVX1 $T=1977360 1108240 0 0 $X=1977358 $Y=1107838
X245 5483 4 2 5477 INVX1 $T=1992540 1128400 1 0 $X=1992538 $Y=1122960
X246 5643 4 2 5596 INVX1 $T=2038740 1098160 0 180 $X=2037420 $Y=1092720
X247 5627 4 2 5597 INVX1 $T=2044020 1098160 1 180 $X=2042700 $Y=1097758
X248 5679 4 2 5664 INVX1 $T=2054580 1027600 1 180 $X=2053260 $Y=1027198
X249 348 4 2 5745 INVX1 $T=2058540 1078000 1 0 $X=2058538 $Y=1072560
X250 347 4 2 5743 INVX1 $T=2058540 1128400 0 0 $X=2058538 $Y=1127998
X251 5662 4 2 5733 INVX1 $T=2059200 987280 1 0 $X=2059198 $Y=981840
X252 5731 4 2 5744 INVX1 $T=2067780 1017520 0 180 $X=2066460 $Y=1012080
X253 374 4 2 5979 INVX1 $T=2135760 1108240 0 0 $X=2135758 $Y=1107838
X254 392 4 2 388 INVX1 $T=2185920 987280 1 0 $X=2185918 $Y=981840
X255 395 4 2 6101 INVX1 $T=2187900 997360 0 180 $X=2186580 $Y=991920
X256 389 4 2 352 INVX1 $T=2211000 1078000 1 0 $X=2210998 $Y=1072560
X257 401 4 2 417 INVX1 $T=2271720 1108240 0 0 $X=2271718 $Y=1107838
X258 411 4 2 6454 INVX1 $T=2298780 1078000 0 0 $X=2298778 $Y=1077598
X259 394 4 2 419 INVX1 $T=2333100 1078000 0 0 $X=2333098 $Y=1077598
X260 6605 4 2 6606 INVX1 $T=2361480 1118320 0 0 $X=2361478 $Y=1117918
X261 6550 4 2 6636 INVX1 $T=2372040 1108240 1 0 $X=2372038 $Y=1102800
X262 6621 4 2 6674 INVX1 $T=2385240 1108240 0 0 $X=2385238 $Y=1107838
X263 420 4 2 6677 INVX1 $T=2390520 1128400 0 0 $X=2390518 $Y=1127998
X264 6675 4 2 6688 INVX1 $T=2393160 1098160 0 0 $X=2393158 $Y=1097758
X265 422 4 2 6704 INVX1 $T=2398440 1118320 0 0 $X=2398438 $Y=1117918
X266 6730 4 2 6741 INVX1 $T=2401080 1108240 1 0 $X=2401078 $Y=1102800
X267 411 4 2 6773 INVX1 $T=2420880 1088080 1 0 $X=2420878 $Y=1082640
X268 7090 4 2 7035 INVX1 $T=2533080 1118320 1 180 $X=2531760 $Y=1117918
X269 1979 47 2 2002 1954 4 AOI21X2 $T=898920 1108240 1 0 $X=898918 $Y=1102800
X270 2222 75 2 2295 2205 4 AOI21X2 $T=995940 1138480 1 0 $X=995938 $Y=1133040
X271 3714 3761 2 3770 3790 4 AOI21X2 $T=1474440 1067920 0 0 $X=1474438 $Y=1067518
X272 3825 3826 2 3789 201 4 AOI21X2 $T=1494240 1017520 0 0 $X=1494238 $Y=1017118
X273 4037 3942 2 3975 4036 4 AOI21X2 $T=1554960 1067920 1 180 $X=1550340 $Y=1067518
X274 4161 4128 2 4194 4222 4 AOI21X2 $T=1604460 1078000 1 180 $X=1599840 $Y=1077598
X275 268 4788 2 4821 4837 4 AOI21X2 $T=1790580 1128400 0 180 $X=1785960 $Y=1122960
X276 5142 5099 2 5133 5123 4 AOI21X2 $T=1878360 1118320 1 180 $X=1873740 $Y=1117918
X277 301 296 2 5204 5205 4 AOI21X2 $T=1896180 987280 1 0 $X=1896178 $Y=981840
X278 5457 5427 2 5477 5456 4 AOI21X2 $T=1984620 1128400 1 0 $X=1984618 $Y=1122960
X279 5758 5731 2 5788 5791 4 AOI21X2 $T=2075700 997360 1 0 $X=2075698 $Y=991920
X280 6968 440 2 6970 6944 4 AOI21X2 $T=2497440 1128400 1 0 $X=2497438 $Y=1122960
X281 2 2038 52 2001 4 NOR2X1 $T=910140 1128400 1 180 $X=908160 $Y=1127998
X282 2 2062 1983 2006 4 NOR2X1 $T=920040 1098160 1 180 $X=918060 $Y=1097758
X283 2 56 57 1983 4 NOR2X1 $T=932580 1108240 0 180 $X=930600 $Y=1102800
X284 2 59 58 2062 4 NOR2X1 $T=937860 1098160 1 180 $X=935880 $Y=1097758
X285 2 61 60 2038 4 NOR2X1 $T=940500 1128400 1 180 $X=938520 $Y=1127998
X286 2 2160 2114 2159 4 NOR2X1 $T=946440 1088080 1 0 $X=946438 $Y=1082640
X287 2 2162 2163 2176 4 NOR2X1 $T=954360 1037680 0 0 $X=954358 $Y=1037278
X288 2 2163 2171 2172 4 NOR2X1 $T=954360 1047760 0 0 $X=954358 $Y=1047358
X289 2 2220 2171 2221 4 NOR2X1 $T=975480 1047760 1 0 $X=975478 $Y=1042320
X290 2 2330 2292 2175 4 NOR2X1 $T=997920 1078000 1 180 $X=995940 $Y=1077598
X291 2 2389 2388 2330 4 NOR2X1 $T=1025640 1078000 0 180 $X=1023660 $Y=1072560
X292 2 2411 81 2222 4 NOR2X1 $T=1029600 1138480 0 180 $X=1027620 $Y=1133040
X293 2 2416 2414 2411 4 NOR2X1 $T=1034220 1128400 0 180 $X=1032240 $Y=1122960
X294 2 2477 2381 2292 4 NOR2X1 $T=1037520 1088080 0 180 $X=1035540 $Y=1082640
X295 2 85 2448 81 4 NOR2X1 $T=1060620 1138480 0 180 $X=1058640 $Y=1133040
X296 2 92 95 111 4 NOR2X1 $T=1114080 997360 0 0 $X=1114078 $Y=996958
X297 2 3110 3104 3144 4 NOR2X1 $T=1252020 1037680 1 0 $X=1252018 $Y=1032240
X298 2 3198 3197 3195 4 NOR2X1 $T=1275120 1057840 1 0 $X=1275118 $Y=1052400
X299 2 3702 3725 3726 4 NOR2X1 $T=1459260 1128400 1 0 $X=1459258 $Y=1122960
X300 2 3635 3731 3729 4 NOR2X1 $T=1463880 1017520 0 180 $X=1461900 $Y=1012080
X301 2 3807 3729 3826 4 NOR2X1 $T=1488300 1027600 1 0 $X=1488298 $Y=1022160
X302 2 202 199 3890 4 NOR2X1 $T=1504140 1128400 0 0 $X=1504138 $Y=1127998
X303 2 4773 4817 4807 4 NOR2X1 $T=1783980 1047760 1 180 $X=1782000 $Y=1047358
X304 2 5648 5689 5642 4 NOR2X1 $T=2051940 1088080 1 180 $X=2049960 $Y=1087678
X305 2 5767 5714 5643 4 NOR2X1 $T=2053260 1098160 1 180 $X=2051280 $Y=1097758
X306 2 5681 5729 5728 4 NOR2X1 $T=2057220 1027600 1 0 $X=2057218 $Y=1022160
X307 2 6185 6149 392 4 NOR2X1 $T=2199120 997360 0 180 $X=2197140 $Y=991920
X308 2 6363 6452 6535 4 NOR2X1 $T=2333760 1128400 1 0 $X=2333758 $Y=1122960
X309 2 6410 6509 6536 4 NOR2X1 $T=2337060 1108240 0 0 $X=2337058 $Y=1107838
X310 2 6536 6535 6550 4 NOR2X1 $T=2339040 1118320 0 0 $X=2339038 $Y=1117918
X311 2 419 6455 6610 4 NOR2X1 $T=2344320 1078000 0 0 $X=2344318 $Y=1077598
X312 2 6610 6635 6612 4 NOR2X1 $T=2372040 1098160 1 0 $X=2372038 $Y=1092720
X313 2 6525 6486 6635 4 NOR2X1 $T=2379960 1098160 1 0 $X=2379958 $Y=1092720
X314 2 6636 6704 6730 4 NOR2X1 $T=2397780 1108240 0 0 $X=2397778 $Y=1107838
X315 2 6775 6702 433 4 NOR2X1 $T=2432100 1118320 0 0 $X=2432098 $Y=1117918
X316 2 438 452 453 4 NOR2X1 $T=2553540 1138480 1 0 $X=2553538 $Y=1133040
X317 1714 1769 4 2 1757 NOR2X2 $T=831600 1118320 1 180 $X=828300 $Y=1117918
X318 1779 38 4 2 1769 NOR2X2 $T=834900 1128400 0 180 $X=831600 $Y=1122960
X319 1777 1715 4 2 1790 NOR2X2 $T=834240 1067920 1 0 $X=834238 $Y=1062480
X320 1778 1685 4 2 1775 NOR2X2 $T=834240 1078000 0 0 $X=834238 $Y=1077598
X321 2558 114 4 2 116 NOR2X2 $T=1136520 1057840 1 0 $X=1136518 $Y=1052400
X322 3595 3557 4 2 3725 NOR2X2 $T=1440120 1118320 0 0 $X=1440118 $Y=1117918
X323 3596 194 4 2 3702 NOR2X2 $T=1441440 1128400 0 0 $X=1441438 $Y=1127998
X324 3793 3788 4 2 3866 NOR2X2 $T=1494900 1118320 0 0 $X=1494898 $Y=1117918
X325 3866 3890 4 2 3927 NOR2X2 $T=1518660 1118320 0 0 $X=1518658 $Y=1117918
X326 4038 3317 4 2 4039 NOR2X2 $T=1558920 1007440 0 180 $X=1555620 $Y=1002000
X327 4039 4008 4 2 4086 NOR2X2 $T=1572120 1017520 1 180 $X=1568820 $Y=1017118
X328 1874 215 4 2 4190 NOR2X2 $T=1598520 1118320 0 0 $X=1598518 $Y=1117918
X329 230 231 4 2 233 NOR2X2 $T=1649340 1037680 0 0 $X=1649338 $Y=1037278
X330 4418 4421 4 2 4419 NOR2X2 $T=1669140 1138480 0 180 $X=1665840 $Y=1133040
X331 4265 4594 4 2 4578 NOR2X2 $T=1721940 1067920 0 180 $X=1718640 $Y=1062480
X332 4802 4772 4 2 4836 NOR2X2 $T=1777380 1088080 0 0 $X=1777378 $Y=1087678
X333 4269 4818 4 2 267 NOR2X2 $T=1788600 997360 1 0 $X=1788598 $Y=991920
X334 4864 267 4 2 4896 NOR2X2 $T=1797180 997360 0 0 $X=1797178 $Y=996958
X335 310 309 4 2 5260 NOR2X2 $T=1912020 1098160 1 180 $X=1908720 $Y=1097758
X336 5260 5291 4 2 5292 NOR2X2 $T=1925880 1108240 0 180 $X=1922580 $Y=1102800
X337 322 323 4 2 5291 NOR2X2 $T=1948320 1108240 1 0 $X=1948318 $Y=1102800
X338 4782 5482 4 2 337 NOR2X2 $T=1990560 987280 0 0 $X=1990558 $Y=986878
X339 5583 5607 4 2 5622 NOR2X2 $T=2024220 1057840 0 0 $X=2024218 $Y=1057438
X340 5594 5592 4 2 5607 NOR2X2 $T=2028180 1067920 0 180 $X=2024880 $Y=1062480
X341 5793 5727 4 2 5758 NOR2X2 $T=2074380 997360 1 180 $X=2071080 $Y=996958
X342 5773 5771 4 2 5681 NOR2X2 $T=2075700 1047760 0 0 $X=2075698 $Y=1047358
X343 5801 5802 4 2 5727 NOR2X2 $T=2090220 1007440 0 0 $X=2090218 $Y=1007038
X344 5830 5832 4 2 5729 NOR2X2 $T=2096820 1027600 0 0 $X=2096818 $Y=1027198
X345 5891 5893 4 2 5793 NOR2X2 $T=2112660 997360 0 0 $X=2112658 $Y=996958
X346 6009 6004 4 2 375 NOR2X2 $T=2147640 997360 0 0 $X=2147638 $Y=996958
X347 6040 6041 4 2 382 NOR2X2 $T=2156220 997360 0 0 $X=2156218 $Y=996958
X348 5891 5893 4 2 5831 OR2XL $T=2103420 997360 1 180 $X=2100780 $Y=996958
X349 1773 1774 1772 4 2 NAND2X2 $T=835560 1037680 0 180 $X=832260 $Y=1032240
X350 1779 38 1792 4 2 NAND2X2 $T=834240 1118320 0 0 $X=834238 $Y=1117918
X351 3264 3229 3245 4 2 NAND2X2 $T=1294920 1078000 0 0 $X=1294918 $Y=1077598
X352 3638 3704 3773 4 2 NAND2X2 $T=1481040 1037680 0 180 $X=1477740 $Y=1032240
X353 3714 3756 3804 4 2 NAND2X2 $T=1488960 1067920 1 180 $X=1485660 $Y=1067518
X354 3986 3366 4060 4 2 NAND2X2 $T=1556940 1027600 1 180 $X=1553640 $Y=1027198
X355 1901 4118 4103 4 2 NAND2X2 $T=1575420 1078000 0 180 $X=1572120 $Y=1072560
X356 1877 211 4130 4 2 NAND2X2 $T=1575420 1108240 1 180 $X=1572120 $Y=1107838
X357 4339 4360 4342 4 2 NAND2X2 $T=1647360 1108240 1 180 $X=1644060 $Y=1107838
X358 4388 4426 4445 4 2 NAND2X2 $T=1671780 1088080 1 0 $X=1671778 $Y=1082640
X359 4494 254 253 4 2 NAND2X2 $T=1692900 1138480 0 180 $X=1689600 $Y=1133040
X360 4493 254 4573 4 2 NAND2X2 $T=1694880 1098160 1 180 $X=1691580 $Y=1097758
X361 4265 4594 4576 4 2 NAND2X2 $T=1718640 1067920 0 0 $X=1718638 $Y=1067518
X362 4546 4623 4621 4 2 NAND2X2 $T=1727880 1108240 0 0 $X=1727878 $Y=1107838
X363 4087 4771 4783 4 2 NAND2X2 $T=1773420 1057840 1 180 $X=1770120 $Y=1057438
X364 5142 5081 5169 4 2 NAND2X2 $T=1886280 1128400 1 0 $X=1886278 $Y=1122960
X365 310 309 5249 4 2 NAND2X2 $T=1912020 1098160 0 180 $X=1908720 $Y=1092720
X366 5457 5410 5453 4 2 NAND2X2 $T=1978680 1138480 1 0 $X=1978678 $Y=1133040
X367 6009 6004 377 4 2 NAND2X2 $T=2147640 1007440 0 0 $X=2147638 $Y=1007038
X368 39 2 1757 1768 4 1850 AOI21X4 $T=840840 1108240 0 0 $X=840838 $Y=1107838
X369 2159 2 63 2173 4 49 AOI21X4 $T=951720 1088080 1 0 $X=951718 $Y=1082640
X370 198 2 3726 3733 4 3734 AOI21X4 $T=1459260 1118320 1 0 $X=1459258 $Y=1112880
X371 3927 2 207 3880 4 4052 AOI21X4 $T=1525920 1118320 0 0 $X=1525918 $Y=1117918
X372 3920 2 3975 3989 4 3990 AOI21X4 $T=1540440 1057840 1 0 $X=1540438 $Y=1052400
X373 4086 2 4050 4069 4 214 AOI21X4 $T=1578060 1017520 0 0 $X=1578058 $Y=1017118
X374 4404 2 4388 4389 4 4390 AOI21X4 $T=1665180 1078000 1 180 $X=1658580 $Y=1077598
X375 4801 2 4803 4789 4 4790 AOI21X4 $T=1782660 1017520 0 180 $X=1776060 $Y=1012080
X376 4896 2 4855 4841 4 274 AOI21X4 $T=1798500 987280 0 0 $X=1798498 $Y=986878
X377 5193 2 5292 5307 4 5310 AOI21X4 $T=1922580 1118320 1 0 $X=1922578 $Y=1112880
X378 5627 2 5622 5639 4 5668 AOI21X4 $T=2032140 1057840 1 0 $X=2032138 $Y=1052400
X379 440 2 7049 7035 4 7000 AOI21X4 $T=2519880 1118320 0 180 $X=2513280 $Y=1112880
X380 31 2 1639 4 1641 AND2X2 $T=794640 1118320 0 0 $X=794638 $Y=1117918
X381 1729 2 1713 4 1756 AND2X2 $T=821700 1118320 0 0 $X=821698 $Y=1117918
X382 1916 2 1927 4 1936 AND2X2 $T=884400 1037680 0 0 $X=884398 $Y=1037278
X383 2006 2 2001 4 2018 AND2X2 $T=904200 1098160 0 0 $X=904198 $Y=1097758
X384 2161 2 2174 4 2097 AND2X2 $T=943140 1017520 0 180 $X=940500 $Y=1012080
X385 2175 2 2197 4 2252 AND2X2 $T=990660 1088080 0 180 $X=988020 $Y=1082640
X386 3229 2 3211 4 3212 AND2X2 $T=1281060 1037680 0 180 $X=1278420 $Y=1032240
X387 3226 2 158 4 3230 AND2X2 $T=1294920 1118320 1 0 $X=1294918 $Y=1112880
X388 159 2 3226 4 3216 AND2X2 $T=1308120 1128400 0 180 $X=1305480 $Y=1122960
X389 173 2 174 4 3478 AND2X2 $T=1365540 1108240 0 0 $X=1365538 $Y=1107838
X390 200 2 205 4 3892 AND2X2 $T=1516020 987280 0 180 $X=1513380 $Y=981840
X391 3942 2 3971 4 4009 AND2X2 $T=1539780 1088080 1 0 $X=1539778 $Y=1082640
X392 3920 2 3957 4 4055 AND2X2 $T=1542420 1067920 1 0 $X=1542418 $Y=1062480
X393 4101 2 4053 4 4169 AND2X2 $T=1580700 1007440 0 0 $X=1580698 $Y=1007038
X394 4127 2 4137 4 4220 AND2X2 $T=1594560 1047760 0 0 $X=1594558 $Y=1047358
X395 4572 2 258 4 4574 AND2X2 $T=1710720 1118320 0 0 $X=1710718 $Y=1117918
X396 4604 2 263 4 4623 AND2X2 $T=1725240 1128400 0 0 $X=1725238 $Y=1127998
X397 5689 2 5648 4 5578 AND2X2 $T=2057880 1088080 0 0 $X=2057878 $Y=1087678
X398 6612 2 6550 4 6640 AND2X2 $T=2374020 1118320 1 0 $X=2374018 $Y=1112880
X399 7002 2 7049 4 6968 AND2X2 $T=2517900 1128400 0 180 $X=2515260 $Y=1122960
X400 7049 2 7090 4 6945 AND2X2 $T=2528460 1118320 1 180 $X=2525820 $Y=1117918
X401 4103 4 4128 2 4156 NAND2X4 $T=1591920 1078000 1 180 $X=1587300 $Y=1077598
X402 215 4 1874 2 4170 NAND2X4 $T=1594560 1118320 1 180 $X=1589940 $Y=1117918
X403 4421 4 4418 2 4413 NAND2X4 $T=1670460 1128400 0 180 $X=1665840 $Y=1122960
X404 254 4 4498 2 4546 NAND2X4 $T=1696860 1108240 0 0 $X=1696858 $Y=1107838
X405 27 28 4 2 1578 OR2X2 $T=762960 1128400 1 0 $X=762958 $Y=1122960
X406 1790 1775 4 2 1771 OR2X2 $T=835560 1067920 1 180 $X=832920 $Y=1067518
X407 1776 1577 4 2 1773 OR2X2 $T=848100 1037680 0 180 $X=845460 $Y=1032240
X408 2286 72 4 2 2209 OR2X2 $T=982740 987280 0 180 $X=980100 $Y=981840
X409 2287 2251 4 2 2161 OR2X2 $T=984060 1007440 0 180 $X=981420 $Y=1002000
X410 2321 67 4 2 2339 OR2X2 $T=1006500 1088080 1 0 $X=1006498 $Y=1082640
X411 2359 2358 4 2 2267 OR2X2 $T=1015080 1017520 1 180 $X=1012440 $Y=1017118
X412 2360 2385 4 2 2268 OR2X2 $T=1025640 1037680 1 180 $X=1023000 $Y=1037278
X413 3199 3152 4 2 3229 OR2X2 $T=1281060 1088080 0 0 $X=1281058 $Y=1087678
X414 164 165 4 2 166 OR2X2 $T=1336500 987280 1 0 $X=1336498 $Y=981840
X415 3606 3582 4 2 3756 OR2X2 $T=1458600 1088080 0 0 $X=1458598 $Y=1087678
X416 1875 4104 4 2 4127 OR2X2 $T=1574760 1047760 0 0 $X=1574758 $Y=1047358
X417 4190 4106 4 2 4221 OR2X2 $T=1598520 1108240 0 0 $X=1598518 $Y=1107838
X418 3929 4787 4 2 4788 OR2X2 $T=1775400 1108240 0 0 $X=1775398 $Y=1107838
X419 4807 4803 4 2 4805 OR2X2 $T=1781340 1037680 1 180 $X=1778700 $Y=1037278
X420 4088 4806 4 2 4808 OR2X2 $T=1779360 1108240 1 0 $X=1779358 $Y=1102800
X421 293 292 4 2 5081 OR2X2 $T=1867140 1128400 0 180 $X=1864500 $Y=1122960
X422 325 326 4 2 5410 OR2X2 $T=1947660 1118320 0 0 $X=1947658 $Y=1117918
X423 5689 5648 4 2 5564 OR2X2 $T=2042040 1088080 1 180 $X=2039400 $Y=1087678
X424 445 446 4 2 7002 OR2X2 $T=2511300 1138480 0 180 $X=2508660 $Y=1133040
X425 28 4 2 27 1591 NAND2XL $T=773520 1128400 0 0 $X=773518 $Y=1127998
X426 35 4 2 34 1639 NAND2XL $T=793980 1138480 0 180 $X=792000 $Y=1133040
X427 1938 4 2 1927 1914 NAND2XL $T=891000 1027600 1 180 $X=889020 $Y=1027198
X428 2172 4 2 2197 2191 NAND2XL $T=964260 1057840 0 0 $X=964258 $Y=1057438
X429 2221 4 2 2197 2219 NAND2XL $T=974160 1057840 1 180 $X=972180 $Y=1057438
X430 2322 4 2 2268 2279 NAND2XL $T=996600 1047760 0 180 $X=994620 $Y=1042320
X431 2323 4 2 2197 2325 NAND2XL $T=1001220 1057840 0 0 $X=1001218 $Y=1057438
X432 97 4 2 2561 2548 NAND2XL $T=1083060 1128400 1 180 $X=1081080 $Y=1127998
X433 97 4 2 2591 2543 NAND2XL $T=1088340 1128400 0 180 $X=1086360 $Y=1122960
X434 3209 4 2 3229 3292 NAND2XL $T=1293600 1088080 0 0 $X=1293598 $Y=1087678
X435 159 4 2 161 3315 NAND2XL $T=1312740 1128400 1 0 $X=1312738 $Y=1122960
X436 4742 4 2 4788 265 NAND2XL $T=1774080 1128400 1 0 $X=1774078 $Y=1122960
X437 4756 4 2 4801 4830 NAND2XL $T=1791240 1017520 0 0 $X=1791238 $Y=1017118
X438 4770 4 2 4808 4910 NAND2XL $T=1807080 1098160 0 0 $X=1807078 $Y=1097758
X439 5080 4 2 5081 5085 NAND2XL $T=1861860 1108240 1 0 $X=1861858 $Y=1102800
X440 298 4 2 5142 5136 NAND2XL $T=1881000 1128400 1 180 $X=1879020 $Y=1127998
X441 5249 4 2 5265 5236 NAND2XL $T=1909380 1088080 0 180 $X=1907400 $Y=1082640
X442 5483 4 2 5457 5428 NAND2XL $T=1986600 1138480 0 180 $X=1984620 $Y=1133040
X443 5628 4 2 5596 5610 NAND2XL $T=2026200 1098160 0 180 $X=2024220 $Y=1092720
X444 6230 4 2 394 6339 NAND2XL $T=2263800 1067920 1 180 $X=2261820 $Y=1067518
X445 394 4 2 383 6338 NAND2XL $T=2270400 1057840 0 180 $X=2268420 $Y=1052400
X446 419 4 2 6455 6609 NAND2XL $T=2346960 1088080 0 0 $X=2346958 $Y=1087678
X447 6563 4 2 6583 6732 NAND2XL $T=2364120 1128400 1 0 $X=2364118 $Y=1122960
X448 6583 4 2 422 6624 NAND2XL $T=2364120 1138480 1 0 $X=2364118 $Y=1133040
X449 394 4 2 6773 6776 NAND2XL $T=2421540 1098160 1 0 $X=2421538 $Y=1092720
X450 454 4 2 456 7211 NAND2XL $T=2560140 1138480 1 0 $X=2560138 $Y=1133040
X451 39 42 4 2 INVX4 $T=853380 1138480 1 0 $X=853378 $Y=1133040
X452 96 100 4 2 INVX4 $T=1129920 1078000 1 0 $X=1129918 $Y=1072560
X453 51 114 4 2 INVX4 $T=1134540 1057840 1 180 $X=1131900 $Y=1057438
X454 163 162 4 2 INVX4 $T=1318020 1078000 1 180 $X=1315380 $Y=1077598
X455 201 204 4 2 INVX4 $T=1504140 997360 0 0 $X=1504138 $Y=996958
X456 4050 4189 4 2 INVX4 $T=1585320 1027600 1 0 $X=1585318 $Y=1022160
X457 5668 5662 4 2 INVX4 $T=2043360 1007440 1 180 $X=2040720 $Y=1007038
X458 31 29 2 1605 1603 4 AOI21X1 $T=776820 1118320 1 0 $X=776818 $Y=1112880
X459 2001 47 2 2007 1977 4 AOI21X1 $T=902880 1118320 0 0 $X=902878 $Y=1117918
X460 2007 2006 2 2034 2017 4 AOI21X1 $T=917400 1088080 0 0 $X=917398 $Y=1087678
X461 2172 2188 2 2190 2192 4 AOI21X1 $T=958980 1047760 0 0 $X=958978 $Y=1047358
X462 2234 2176 2 2193 2194 4 AOI21X1 $T=964260 1078000 0 180 $X=961620 $Y=1072560
X463 2217 2209 2 2207 2195 4 AOI21X1 $T=970860 997360 1 180 $X=968220 $Y=996958
X464 2161 2249 2 2217 2218 4 AOI21X1 $T=982740 1017520 1 180 $X=980100 $Y=1017118
X465 2175 2188 2 2234 2253 4 AOI21X1 $T=989340 1078000 0 180 $X=986700 $Y=1072560
X466 2278 2188 2 2272 2288 4 AOI21X1 $T=993300 1088080 0 0 $X=993298 $Y=1087678
X467 2323 2188 2 2329 2320 4 AOI21X1 $T=1002540 1057840 1 0 $X=1002538 $Y=1052400
X468 95 92 2 111 112 4 AOI21X1 $T=1117380 987280 0 0 $X=1117378 $Y=986878
X469 3015 2796 2 3058 156 4 AOI21X1 $T=1236180 997360 0 0 $X=1236178 $Y=996958
X470 3091 3192 2 3195 3196 4 AOI21X1 $T=1271820 1017520 0 0 $X=1271818 $Y=1017118
X471 3756 3801 2 3761 3809 4 AOI21X1 $T=1485660 1088080 0 0 $X=1485658 $Y=1087678
X472 5081 5084 2 5099 5139 4 AOI21X1 $T=1875720 1108240 1 0 $X=1875718 $Y=1102800
X473 5410 5425 2 5427 5426 4 AOI21X1 $T=1968780 1128400 1 0 $X=1968778 $Y=1122960
X474 5662 5682 2 5684 345 4 AOI21X1 $T=2047320 1007440 0 0 $X=2047318 $Y=1007038
X475 5728 5662 2 5731 5712 4 AOI21X1 $T=2057880 997360 1 0 $X=2057878 $Y=991920
X476 388 381 2 6101 390 4 AOI21X1 $T=2179320 987280 1 0 $X=2179318 $Y=981840
X477 6621 6612 2 6611 6605 4 AOI21X1 $T=2367420 1108240 0 180 $X=2364780 $Y=1102800
X478 6640 420 2 6606 6703 4 AOI21X1 $T=2379300 1118320 0 0 $X=2379298 $Y=1117918
X479 1714 1792 4 1713 2 1768 OAI21X2 $T=832260 1108240 1 180 $X=826980 $Y=1107838
X480 1771 1850 4 1803 2 1848 OAI21X2 $T=852060 1057840 1 0 $X=852058 $Y=1052400
X481 3804 3734 4 3790 2 3825 OAI21X2 $T=1493580 1067920 0 0 $X=1493578 $Y=1067518
X482 3807 3839 4 3773 2 3840 OAI21X2 $T=1498860 1027600 1 180 $X=1493580 $Y=1027198
X483 3866 203 4 3823 2 3880 OAI21X2 $T=1508760 1118320 1 180 $X=1503480 $Y=1117918
X484 4060 4039 4 4053 2 4069 OAI21X2 $T=1562880 1017520 1 180 $X=1557600 $Y=1017118
X485 4106 4170 4 4130 2 4161 OAI21X2 $T=1594560 1108240 1 180 $X=1589280 $Y=1107838
X486 4008 4189 4 4060 2 4198 OAI21X2 $T=1599840 1017520 1 180 $X=1594560 $Y=1017118
X487 217 4221 4 4236 2 4253 OAI21X2 $T=1615680 1098160 1 180 $X=1610400 $Y=1097758
X488 241 4419 4 4413 2 4473 OAI21X2 $T=1678380 1118320 1 180 $X=1673100 $Y=1117918
X489 241 4438 4 4446 2 4466 OAI21X2 $T=1681020 1088080 1 180 $X=1675740 $Y=1087678
X490 5291 5249 4 5303 2 5307 OAI21X2 $T=1921920 1098160 1 0 $X=1921918 $Y=1092720
X491 5679 5729 4 5742 2 5731 OAI21X2 $T=2073060 1027600 1 0 $X=2073058 $Y=1022160
X492 1772 1848 1875 4 2 XNOR2X4 $T=849420 1047760 0 0 $X=849418 $Y=1047358
X493 2279 2260 78 4 2 XNOR2X4 $T=991320 1108240 0 0 $X=991318 $Y=1107838
X494 3803 3840 3986 4 2 XNOR2X4 $T=1508100 1027600 0 0 $X=1508098 $Y=1027198
X495 4055 4036 4087 4 2 XNOR2X4 $T=1560240 1067920 1 0 $X=1560238 $Y=1062480
X496 4156 4253 4326 4 2 XNOR2X4 $T=1611720 1088080 1 0 $X=1611718 $Y=1082640
X497 4548 4444 4498 4 2 XNOR2X4 $T=1704780 1067920 1 180 $X=1693560 $Y=1067518
X498 4830 4805 269 4 2 XNOR2X4 $T=1787940 1037680 0 0 $X=1787938 $Y=1037278
X499 5667 5662 5503 4 2 XNOR2X4 $T=2049960 997360 1 180 $X=2038740 $Y=996958
X500 5950 5947 370 4 2 XNOR2X4 $T=2129820 987280 0 180 $X=2118600 $Y=981840
X501 1769 4 42 1792 2 1861 OAI21X4 $T=853380 1128400 1 0 $X=853378 $Y=1122960
X502 4052 4 4051 3990 2 4050 OAI21X4 $T=1559580 1057840 0 180 $X=1552320 $Y=1052400
X503 4190 4 217 4170 2 4249 OAI21X4 $T=1613040 1108240 1 180 $X=1605780 $Y=1107838
X504 4239 4 217 4222 2 4235 OAI21X4 $T=1613700 1078000 0 180 $X=1606440 $Y=1072560
X505 4413 4 4382 4342 2 4404 OAI21X4 $T=1667160 1108240 1 180 $X=1659900 $Y=1107838
X506 241 4 4445 4390 2 4444 OAI21X4 $T=1678380 1078000 0 180 $X=1671120 $Y=1072560
X507 267 4 4790 266 2 4841 OAI21X4 $T=1793220 987280 1 180 $X=1785960 $Y=986878
X508 4853 4 4852 4836 2 4855 OAI21X4 $T=1798500 1088080 1 180 $X=1791240 $Y=1087678
X509 302 4 5169 5123 2 5193 OAI21X4 $T=1885620 1118320 1 0 $X=1885618 $Y=1112880
X510 5453 4 5310 5456 2 333 OAI21X4 $T=1974720 1128400 1 0 $X=1974718 $Y=1122960
X511 338 4 5641 339 2 5627 OAI21X4 $T=2036760 1128400 0 0 $X=2036758 $Y=1127998
X512 5733 4 5772 5791 2 5880 OAI21X4 $T=2074380 987280 1 0 $X=2074378 $Y=981840
X513 375 4 369 377 2 5947 OAI21X4 $T=2136420 987280 1 0 $X=2136418 $Y=981840
X514 1601 1603 2 4 1715 XOR2X2 $T=775500 1098160 1 0 $X=775498 $Y=1092720
X515 1641 29 2 4 1685 XOR2X2 $T=792660 1108240 0 0 $X=792658 $Y=1107838
X516 1958 1954 2 4 1698 XOR2X2 $T=894300 1108240 0 180 $X=887700 $Y=1102800
X517 3808 3809 2 4 3909 XOR2X2 $T=1486980 1078000 0 0 $X=1486978 $Y=1077598
X518 3867 3839 2 4 3908 XOR2X2 $T=1501500 1047760 0 0 $X=1501498 $Y=1047358
X519 3892 204 2 4 4038 XOR2X2 $T=1512060 997360 0 0 $X=1512058 $Y=996958
X520 3907 3921 2 4 3929 XOR2X2 $T=1519320 1108240 0 0 $X=1519318 $Y=1107838
X521 4223 4189 2 4 4267 XOR2X2 $T=1603800 1027600 1 0 $X=1603798 $Y=1022160
X522 4910 4837 2 4 275 XOR2X2 $T=1804440 1128400 1 0 $X=1804438 $Y=1122960
X523 6945 440 2 4 6934 XOR2X2 $T=2490180 1118320 0 180 $X=2483580 $Y=1112880
X524 7001 7000 2 4 6969 XOR2X2 $T=2504700 1098160 1 180 $X=2498100 $Y=1097758
X525 2205 4 2188 2 INVX2 $T=967560 1088080 0 0 $X=967558 $Y=1087678
X526 2114 4 2197 2 INVX2 $T=972180 1088080 1 0 $X=972178 $Y=1082640
X527 3293 4 3463 2 INVX2 $T=1314720 1067920 1 0 $X=1314718 $Y=1062480
X528 3759 4 3761 2 INVX2 $T=1471800 1088080 0 0 $X=1471798 $Y=1087678
X529 3734 4 3801 2 INVX2 $T=1495560 1098160 1 0 $X=1495558 $Y=1092720
X530 3971 4 3975 2 INVX2 $T=1537800 1078000 0 0 $X=1537798 $Y=1077598
X531 4381 4 4389 2 INVX2 $T=1652640 1078000 0 0 $X=1652638 $Y=1077598
X532 4426 4 4438 2 INVX2 $T=1671120 1088080 0 0 $X=1671118 $Y=1087678
X533 4783 4 4803 2 INVX2 $T=1775400 1057840 1 0 $X=1775398 $Y=1052400
X534 2175 2 4 2171 INVXL $T=958320 1057840 0 180 $X=957000 $Y=1052400
X535 2281 2 4 2272 INVXL $T=991980 1088080 1 180 $X=990660 $Y=1087678
X536 2292 2 4 2278 INVXL $T=995280 1088080 0 180 $X=993960 $Y=1082640
X537 2835 2 4 131 INVXL $T=1183380 987280 0 0 $X=1183378 $Y=986878
X538 219 2 4 4403 INVXL $T=1664520 1047760 1 180 $X=1663200 $Y=1047358
X539 5099 2 4 5080 INVXL $T=1866480 1108240 0 180 $X=1865160 $Y=1102800
X540 300 2 4 5204 INVXL $T=1906740 987280 1 0 $X=1906738 $Y=981840
X541 5260 2 4 5265 INVXL $T=1917300 1088080 0 180 $X=1915980 $Y=1082640
X542 394 2 4 6030 INVXL $T=2187900 1078000 1 180 $X=2186580 $Y=1077598
X543 6535 2 4 6583 INVXL $T=2340360 1128400 1 0 $X=2340358 $Y=1122960
X544 6635 2 4 6687 INVXL $T=2385240 1088080 0 0 $X=2385238 $Y=1087678
X545 1578 31 29 2 1567 1566 4 AOI31X1 $T=766920 1118320 0 180 $X=763620 $Y=1112880
X546 2282 2280 2 4 73 XNOR2X2 $T=995280 1057840 1 180 $X=988020 $Y=1057438
X547 2344 2341 2 4 77 XNOR2X2 $T=1010460 1098160 1 180 $X=1003200 $Y=1097758
X548 3747 3743 2 4 199 XNOR2X2 $T=1467840 1128400 0 0 $X=1467838 $Y=1127998
X549 4411 4466 2 4 4493 XNOR2X2 $T=1683660 1088080 1 0 $X=1683658 $Y=1082640
X550 4481 4473 2 4 4494 XNOR2X2 $T=1686300 1118320 0 0 $X=1686298 $Y=1117918
X551 270 4863 2 4 272 XNOR2X2 $T=1798500 987280 1 0 $X=1798498 $Y=981840
X552 6732 6691 2 4 429 XNOR2X2 $T=2404380 1128400 0 0 $X=2404378 $Y=1127998
X553 26 1566 4 2 1577 XOR2X1 $T=761640 1108240 1 0 $X=761638 $Y=1102800
X554 1938 1936 4 2 1777 XOR2X1 $T=888360 1047760 1 180 $X=883080 $Y=1047358
X555 1927 1916 4 2 1778 XOR2X1 $T=888360 1067920 0 180 $X=883080 $Y=1062480
X556 1976 1977 4 2 1779 XOR2X1 $T=898920 1118320 0 180 $X=893640 $Y=1112880
X557 2097 2158 4 2 65 XOR2X1 $T=948420 1067920 1 0 $X=948418 $Y=1062480
X558 2259 2250 4 2 71 XOR2X1 $T=987360 1108240 0 180 $X=982080 $Y=1102800
X559 99 98 4 2 2573 XOR2X1 $T=1092300 1017520 1 180 $X=1087020 $Y=1017118
X560 119 120 4 2 2676 XOR2X1 $T=1146420 1088080 1 180 $X=1141140 $Y=1087678
X561 118 119 4 2 2726 XOR2X1 $T=1143780 1017520 1 0 $X=1143778 $Y=1012080
X562 2810 129 4 2 2797 XOR2X1 $T=1172160 1118320 1 180 $X=1166880 $Y=1117918
X563 108 104 4 2 2827 XOR2X1 $T=1174800 1047760 0 0 $X=1174798 $Y=1047358
X564 2888 89 4 2 142 XOR2X1 $T=1197240 1037680 1 0 $X=1197238 $Y=1032240
X565 142 2951 4 2 3015 XOR2X1 $T=1209120 1007440 1 0 $X=1209118 $Y=1002000
X566 141 2948 4 2 3105 XOR2X1 $T=1209120 1098160 1 0 $X=1209118 $Y=1092720
X567 2931 2849 4 2 3049 XOR2X1 $T=1209780 1067920 1 0 $X=1209778 $Y=1062480
X568 2972 143 4 2 2951 XOR2X1 $T=1216380 997360 0 180 $X=1211100 $Y=991920
X569 3051 3049 4 2 3117 XOR2X1 $T=1238820 1067920 1 0 $X=1238818 $Y=1062480
X570 149 3117 4 2 3198 XOR2X1 $T=1247400 1057840 0 0 $X=1247398 $Y=1057438
X571 3197 3198 4 2 3263 XOR2X1 $T=1274460 1067920 1 0 $X=1274458 $Y=1062480
X572 174 173 4 2 3500 XOR2X1 $T=1364880 1118320 0 0 $X=1364878 $Y=1117918
X573 4804 4817 4 2 271 XOR2X1 $T=1796520 1057840 0 0 $X=1796518 $Y=1057438
X574 5136 5139 4 2 5152 XOR2X1 $T=1877040 1088080 0 0 $X=1877038 $Y=1087678
X575 5236 5235 4 2 5202 XOR2X1 $T=1902120 1078000 1 180 $X=1896840 $Y=1077598
X576 306 5205 4 2 307 XOR2X1 $T=1898160 987280 0 0 $X=1898158 $Y=986878
X577 5428 5426 4 2 5399 XOR2X1 $T=1971420 1138480 0 180 $X=1966140 $Y=1133040
X578 5441 5425 4 2 5324 XOR2X1 $T=1974060 1108240 1 180 $X=1968780 $Y=1107838
X579 5503 5492 4 2 4818 XOR2X1 $T=1999800 997360 1 180 $X=1994520 $Y=996958
X580 5610 5597 4 2 4787 XOR2X1 $T=2028840 1098160 1 180 $X=2023560 $Y=1097758
X581 5713 5712 4 2 341 XOR2X1 $T=2052600 987280 1 180 $X=2047320 $Y=986878
X582 6259 6230 4 2 6206 XOR2X1 $T=2238060 1057840 1 180 $X=2232780 $Y=1057438
X583 383 394 4 2 6259 XOR2X1 $T=2248620 1057840 1 180 $X=2243340 $Y=1057438
X584 1916 2 1914 1776 4 NOR2BX1 $T=879120 1027600 1 180 $X=876480 $Y=1027198
X585 2001 2 1983 1979 4 NOR2BX1 $T=901560 1098160 0 180 $X=898920 $Y=1092720
X586 3823 2 3866 3907 4 NOR2BX1 $T=1505460 1108240 0 0 $X=1505458 $Y=1107838
X587 212 2 213 4172 4 NOR2BX1 $T=1593240 1088080 0 0 $X=1593238 $Y=1087678
X588 4413 2 4419 240 4 NOR2BX1 $T=1674420 1138480 1 0 $X=1674418 $Y=1133040
X589 4808 2 4742 4802 4 NOR2BX1 $T=1781340 1098160 0 180 $X=1778700 $Y=1092720
X590 5728 2 5727 5682 4 NOR2BX1 $T=2059200 1007440 1 180 $X=2056560 $Y=1007038
X591 411 2 394 6775 4 NOR2BX1 $T=2420220 1118320 1 0 $X=2420218 $Y=1112880
X592 2476 2449 2441 2358 2 4 2385 ADDFX2 $T=1052700 1017520 1 180 $X=1038840 $Y=1017118
X593 2492 84 83 2286 2 4 2287 ADDFX2 $T=1061940 987280 0 180 $X=1048080 $Y=981840
X594 2506 2489 2478 2381 2 4 2416 ADDFX2 $T=1061940 1098160 1 180 $X=1048080 $Y=1097758
X595 2542 86 2488 2251 2 4 2359 ADDFX2 $T=1065240 1007440 0 180 $X=1051380 $Y=1002000
X596 2540 2508 2490 2360 2 4 2389 ADDFX2 $T=1067220 1037680 1 180 $X=1053360 $Y=1037278
X597 2529 2510 2493 2388 2 4 2477 ADDFX2 $T=1067880 1067920 1 180 $X=1054020 $Y=1067518
X598 2528 2519 2504 2492 2 4 2488 ADDFX2 $T=1070520 997360 0 180 $X=1056660 $Y=991920
X599 91 51 88 2504 2 4 2449 ADDFX2 $T=1078440 1017520 1 180 $X=1064580 $Y=1017118
X600 2566 2547 2532 2478 2 4 2527 ADDFX2 $T=1083720 1098160 1 180 $X=1069860 $Y=1097758
X601 2560 93 2527 2414 2 4 2448 ADDFX2 $T=1083720 1118320 0 180 $X=1069860 $Y=1112880
X602 2576 2563 2550 2542 2 4 2441 ADDFX2 $T=1089660 1007440 1 180 $X=1075800 $Y=1007038
X603 2558 96 2556 2510 2 4 2541 ADDFX2 $T=1090320 1067920 1 180 $X=1076460 $Y=1067518
X604 2586 2573 2557 2476 2 4 2540 ADDFX2 $T=1090980 1037680 0 180 $X=1077120 $Y=1032240
X605 2604 2574 2541 2493 2 4 2506 ADDFX2 $T=1090980 1078000 1 180 $X=1077120 $Y=1077598
X606 100 87 2558 2550 2 4 2508 ADDFX2 $T=1091640 1037680 1 180 $X=1077780 $Y=1037278
X607 96 106 102 2547 2 4 2561 ADDFX2 $T=1106160 1098160 1 180 $X=1092300 $Y=1097758
X608 106 107 103 2574 2 4 2566 ADDFX2 $T=1107480 1088080 1 180 $X=1093620 $Y=1087678
X609 110 108 104 2596 2 4 2591 ADDFX2 $T=1107480 1108240 1 180 $X=1093620 $Y=1107838
X610 2626 2625 2606 2490 2 4 2529 ADDFX2 $T=1109460 1057840 0 180 $X=1095600 $Y=1052400
X611 115 99 102 2626 2 4 2604 ADDFX2 $T=1112760 1067920 0 180 $X=1098900 $Y=1062480
X612 88 92 109 2557 2 4 2606 ADDFX2 $T=1116720 1037680 0 180 $X=1102860 $Y=1032240
X613 2676 109 2596 2489 2 4 2532 ADDFX2 $T=1128600 1098160 1 180 $X=1114740 $Y=1097758
X614 168 3436 3452 3453 2 4 3462 ADDFX2 $T=1353000 1078000 1 0 $X=1352998 $Y=1072560
X615 171 172 3478 3436 2 4 3529 ADDFX2 $T=1361580 1088080 0 0 $X=1361578 $Y=1087678
X616 3460 176 178 179 2 4 3590 ADDFX2 $T=1364880 1007440 1 0 $X=1364878 $Y=1002000
X617 168 170 3504 3505 2 4 3527 ADDFX2 $T=1380060 1047760 1 0 $X=1380058 $Y=1042320
X618 3500 171 177 3515 2 4 3520 ADDFX2 $T=1381380 1067920 0 0 $X=1381378 $Y=1067518
X619 180 176 3517 3521 2 4 3578 ADDFX2 $T=1382700 1088080 1 0 $X=1382698 $Y=1082640
X620 168 183 177 3517 2 4 3522 ADDFX2 $T=1383360 1098160 1 0 $X=1383358 $Y=1092720
X621 3478 172 183 3518 2 4 3504 ADDFX2 $T=1387320 1078000 1 0 $X=1387318 $Y=1072560
X622 180 3518 187 3555 2 4 3523 ADDFX2 $T=1389300 997360 0 0 $X=1389298 $Y=996958
X623 3508 3522 3532 3557 2 4 3596 ADDFX2 $T=1390620 1128400 1 0 $X=1390618 $Y=1122960
X624 3519 3529 187 3558 2 4 3532 ADDFX2 $T=1393260 1108240 1 0 $X=1393258 $Y=1102800
X625 180 3461 187 3567 2 4 3581 ADDFX2 $T=1397220 1047760 0 0 $X=1397218 $Y=1047358
X626 3521 3581 3593 3604 2 4 3606 ADDFX2 $T=1409760 1067920 0 0 $X=1409758 $Y=1067518
X627 189 162 3555 192 2 4 3663 ADDFX2 $T=1411080 987280 0 0 $X=1411078 $Y=986878
X628 190 3590 3526 193 2 4 3609 ADDFX2 $T=1411740 1007440 0 0 $X=1411738 $Y=1007038
X629 3622 3663 3609 196 2 4 3724 ADDFX2 $T=1446060 1007440 1 0 $X=1446058 $Y=1002000
X630 361 362 5881 5890 2 4 5715 ADDFX2 $T=2093520 1118320 0 0 $X=2093518 $Y=1117918
X631 5909 5905 364 5832 2 4 5773 ADDFX2 $T=2113980 1067920 1 180 $X=2100120 $Y=1067518
X632 5890 367 5894 5771 2 4 5594 ADDFX2 $T=2117280 1098160 0 180 $X=2103420 $Y=1092720
X633 365 366 368 5919 2 4 5881 ADDFX2 $T=2105400 1128400 1 0 $X=2105398 $Y=1122960
X634 5948 5921 5907 5893 2 4 5801 ADDFX2 $T=2122560 1017520 1 180 $X=2108700 $Y=1017118
X635 371 5932 5918 5802 2 4 5830 ADDFX2 $T=2124540 1027600 1 180 $X=2110680 $Y=1027198
X636 348 353 372 5951 2 4 5905 ADDFX2 $T=2140380 1078000 0 180 $X=2126520 $Y=1072560
X637 5979 5919 373 5909 2 4 5894 ADDFX2 $T=2141040 1118320 1 180 $X=2127180 $Y=1117918
X638 6054 376 5951 5948 2 4 5918 ADDFX2 $T=2144340 1067920 1 180 $X=2130480 $Y=1067518
X639 378 348 383 6027 2 4 5932 ADDFX2 $T=2145000 1027600 1 0 $X=2144998 $Y=1022160
X640 358 380 374 6031 2 4 6044 ADDFX2 $T=2147640 1098160 0 0 $X=2147638 $Y=1097758
X641 6044 383 6027 6012 2 4 5907 ADDFX2 $T=2161500 1037680 0 180 $X=2147640 $Y=1032240
X642 379 365 384 6045 2 4 6054 ADDFX2 $T=2149620 1118320 0 0 $X=2149618 $Y=1117918
X643 6045 386 6030 6007 2 4 5921 ADDFX2 $T=2164140 1088080 0 180 $X=2150280 $Y=1082640
X644 6083 387 6031 6002 2 4 6026 ADDFX2 $T=2164140 1108240 1 180 $X=2150280 $Y=1107838
X645 358 391 389 6086 2 4 6083 ADDFX2 $T=2188560 1108240 1 180 $X=2174700 $Y=1107838
X646 398 353 396 6125 2 4 6029 ADDFX2 $T=2200440 1057840 0 180 $X=2186580 $Y=1052400
X647 6125 6139 6113 6126 2 4 6057 ADDFX2 $T=2200440 1067920 0 180 $X=2186580 $Y=1062480
X648 6205 6215 6206 6203 2 4 6184 ADDFX2 $T=2223540 1027600 1 180 $X=2209680 $Y=1027198
X649 353 401 348 6205 2 4 6139 ADDFX2 $T=2224200 1057840 1 180 $X=2210340 $Y=1057438
X650 365 407 403 6230 2 4 6135 ADDFX2 $T=2234100 1098160 0 180 $X=2220240 $Y=1092720
X651 6263 6228 6247 405 2 4 6192 ADDFX2 $T=2240040 1037680 1 180 $X=2226180 $Y=1037278
X652 389 368 410 408 2 4 404 ADDFX2 $T=2242680 987280 1 180 $X=2228820 $Y=986878
X653 368 414 410 409 2 4 406 ADDFX2 $T=2242680 1007440 1 180 $X=2228820 $Y=1007038
X654 396 348 6261 413 2 4 412 ADDFX2 $T=2247300 1007440 0 180 $X=2233440 $Y=1002000
X655 383 401 416 6363 2 4 418 ADDFX2 $T=2263800 1138480 1 0 $X=2263798 $Y=1133040
X656 398 394 417 6410 2 4 6452 ADDFX2 $T=2282280 1108240 1 0 $X=2282278 $Y=1102800
X657 401 403 6454 6455 2 4 6486 ADDFX2 $T=2292840 1088080 0 0 $X=2292838 $Y=1087678
X658 396 411 419 6525 2 4 6509 ADDFX2 $T=2319900 1098160 1 0 $X=2319898 $Y=1092720
X659 2004 2003 4 2 1938 XNOR2X1 $T=904200 997360 0 180 $X=898920 $Y=991920
X660 2233 2231 4 2 68 XNOR2X1 $T=978780 1067920 1 180 $X=973500 $Y=1067518
X661 2365 80 4 2 79 XNOR2X1 $T=1016400 1138480 0 180 $X=1011120 $Y=1133040
X662 112 91 4 2 2795 XNOR2X1 $T=1134540 987280 0 0 $X=1134538 $Y=986878
X663 107 104 4 2 118 XNOR2X1 $T=1150380 1027600 1 180 $X=1145100 $Y=1027198
X664 120 103 4 2 126 XNOR2X1 $T=1168200 1078000 1 180 $X=1162920 $Y=1077598
X665 120 102 4 2 2810 XNOR2X1 $T=1166880 1108240 0 0 $X=1166878 $Y=1107838
X666 2827 110 4 2 2786 XNOR2X1 $T=1180080 1037680 1 180 $X=1174800 $Y=1037278
X667 2835 122 4 2 134 XNOR2X1 $T=1180080 987280 1 0 $X=1180078 $Y=981840
X668 95 110 4 2 2948 XNOR2X1 $T=1191960 1098160 1 0 $X=1191958 $Y=1092720
X669 2931 102 4 2 138 XNOR2X1 $T=1202520 1017520 1 180 $X=1197240 $Y=1017118
X670 140 137 4 2 2888 XNOR2X1 $T=1202520 1128400 1 180 $X=1197240 $Y=1127998
X671 96 137 4 2 2931 XNOR2X1 $T=1199880 1067920 1 0 $X=1199878 $Y=1062480
X672 137 154 4 2 3118 XNOR2X1 $T=1245420 1128400 0 0 $X=1245418 $Y=1127998
X673 3263 3273 4 2 3293 XNOR2X1 $T=1296240 1067920 1 0 $X=1296238 $Y=1062480
X674 3792 3801 4 2 3793 XNOR2X1 $T=1485000 1108240 1 0 $X=1484998 $Y=1102800
X675 213 212 4 2 4118 XNOR2X1 $T=1582680 1088080 1 180 $X=1577400 $Y=1087678
X676 5085 5084 4 2 5065 XNOR2X1 $T=1866480 1098160 0 180 $X=1861200 $Y=1092720
X677 5348 5300 4 2 5337 XNOR2X1 $T=1943700 1078000 1 180 $X=1938420 $Y=1077598
X678 5563 5580 4 2 4806 XNOR2X1 $T=2018280 1098160 1 180 $X=2013000 $Y=1097758
X679 6041 6040 4 2 5950 XNOR2X1 $T=2159520 987280 0 180 $X=2154240 $Y=981840
X680 6673 6740 4 2 428 XNOR2X1 $T=2405700 1108240 0 0 $X=2405698 $Y=1107838
X681 6742 6660 4 2 427 XNOR2X1 $T=2408340 1088080 0 0 $X=2408338 $Y=1087678
X682 6834 6774 4 2 438 XNOR2X1 $T=2447280 1128400 1 0 $X=2447278 $Y=1122960
X683 7211 455 4 2 7149 XNOR2X1 $T=2562780 1128400 0 180 $X=2557500 $Y=1122960
X684 87 2519 89 2 4 90 ADDHXL $T=1066560 987280 0 0 $X=1066558 $Y=986878
X685 92 2563 95 2 4 2528 ADDHXL $T=1088340 997360 1 180 $X=1081080 $Y=996958
X686 107 2625 105 2 4 2586 ADDHXL $T=1105500 1047760 1 180 $X=1098240 $Y=1047358
X687 4505 4545 250 2 4 4547 ADDHXL $T=1696200 1017520 1 0 $X=1696198 $Y=1012080
X688 257 4544 245 2 4 4505 ADDHXL $T=1704120 997360 0 180 $X=1696860 $Y=991920
X689 291 4991 4977 2 4 5020 ADDHXL $T=1855260 1128400 0 180 $X=1848000 $Y=1122960
X690 5020 4993 5002 2 4 5106 ADDHXL $T=1850640 1098160 0 0 $X=1850638 $Y=1097758
X691 5106 5087 4992 2 4 5120 ADDHXL $T=1866480 1078000 1 0 $X=1866478 $Y=1072560
X692 5120 5151 5016 2 4 5191 ADDHXL $T=1877700 1067920 1 0 $X=1877698 $Y=1062480
X693 5191 5234 5162 2 4 5262 ADDHXL $T=1896180 1067920 1 0 $X=1896178 $Y=1062480
X694 5273 5279 5264 2 4 5288 ADDHXL $T=1915320 1078000 1 0 $X=1915318 $Y=1072560
X695 5288 5289 312 2 4 317 ADDHXL $T=1916640 1128400 0 0 $X=1916638 $Y=1127998
X696 5262 5278 5274 2 4 5273 ADDHXL $T=1923900 1067920 0 180 $X=1916640 $Y=1062480
X697 43 44 45 4 2 1927 XOR3X2 $T=881100 987280 1 0 $X=881098 $Y=981840
X698 97 2561 2591 4 2 101 XOR3X2 $T=1104180 1128400 1 180 $X=1092300 $Y=1127998
X699 2726 125 2797 4 2 2799 XOR3X2 $T=1155000 1047760 1 0 $X=1154998 $Y=1042320
X700 2989 147 2799 4 2 3110 XOR3X2 $T=1223640 1047760 1 0 $X=1223638 $Y=1042320
X701 88 3046 148 4 2 3090 XOR3X2 $T=1225620 1088080 0 0 $X=1225618 $Y=1087678
X702 3090 2971 152 4 2 3152 XOR3X2 $T=1247400 1088080 0 0 $X=1247398 $Y=1087678
X703 3315 158 3226 4 2 3295 XOR3X2 $T=1314060 1128400 1 180 $X=1302180 $Y=1127998
X704 179 186 182 4 2 191 XOR3X2 $T=1391280 987280 1 0 $X=1391278 $Y=981840
X705 3663 3622 3609 4 2 3731 XOR3X2 $T=1445400 1007440 0 0 $X=1445398 $Y=1007038
X706 5613 5594 5592 4 2 4771 XOR3X2 $T=2030820 1078000 0 180 $X=2018940 $Y=1072560
X707 2221 2188 2 2226 4 2225 AOI21XL $T=973500 1047760 0 0 $X=973498 $Y=1047358
X708 1605 1578 1591 4 1567 2 OAI2BB1X1 $T=774840 1118320 1 180 $X=771540 $Y=1117918
X709 2032 2007 2019 4 2002 2 OAI2BB1X1 $T=910800 1108240 0 180 $X=907500 $Y=1102800
X710 63 2252 2253 4 2260 2 OAI2BB1X1 $T=982740 1088080 1 0 $X=982738 $Y=1082640
X711 2267 2294 2283 4 2249 2 OAI2BB1X1 $T=995940 1017520 1 180 $X=992640 $Y=1017118
X712 2268 2234 2322 4 2329 2 OAI2BB1X1 $T=1001880 1047760 1 0 $X=1001878 $Y=1042320
X713 115 96 2710 4 117 2 OAI2BB1X1 $T=1146420 1067920 0 180 $X=1143120 $Y=1062480
X714 2714 2784 2776 4 2796 2 OAI2BB1X1 $T=1158960 1027600 1 0 $X=1158958 $Y=1022160
X715 2797 2726 125 4 2776 2 OAI2BB1X1 $T=1162260 1037680 0 180 $X=1158960 $Y=1032240
X716 2795 2786 123 4 2823 2 OAI2BB1X1 $T=1172820 997360 1 0 $X=1172818 $Y=991920
X717 141 2849 2947 4 2971 2 OAI2BB1X1 $T=1208460 1078000 1 0 $X=1208458 $Y=1072560
X718 142 143 2972 4 144 2 OAI2BB1X1 $T=1211100 987280 0 0 $X=1211098 $Y=986878
X719 148 3046 3045 4 3051 2 OAI2BB1X1 $T=1232220 1078000 1 0 $X=1232218 $Y=1072560
X720 3049 149 3069 4 3104 2 OAI2BB1X1 $T=1237500 1057840 0 0 $X=1237498 $Y=1057438
X721 3105 3118 155 4 3140 2 OAI2BB1X1 $T=1248060 1108240 0 0 $X=1248058 $Y=1107838
X722 3090 152 3142 4 3197 2 OAI2BB1X1 $T=1252020 1088080 1 0 $X=1252018 $Y=1082640
X723 3242 3211 3141 4 3241 2 OAI2BB1X1 $T=1291620 1037680 0 180 $X=1288320 $Y=1032240
X724 206 207 203 4 3921 2 OAI2BB1X1 $T=1519980 1128400 0 0 $X=1519978 $Y=1127998
X725 7035 7002 7015 4 6970 2 OAI2BB1X1 $T=2508660 1118320 1 180 $X=2505360 $Y=1117918
X726 2163 4 2161 2 2220 NAND2BXL $T=974820 1037680 0 180 $X=972180 $Y=1032240
X727 2330 4 2335 2 2344 NAND2BXL $T=1010460 1078000 0 0 $X=1010458 $Y=1077598
X728 5291 4 5303 2 5348 NAND2BXL $T=1941060 1098160 1 0 $X=1941058 $Y=1092720
X729 6610 4 6609 2 6660 NAND2BXL $T=2368740 1088080 0 0 $X=2368738 $Y=1087678
X730 6635 4 6593 2 6673 NAND2BXL $T=2384580 1098160 0 0 $X=2384578 $Y=1097758
X731 169 170 175 3461 2 4 3452 ADDFHX1 $T=1353660 1047760 0 0 $X=1353658 $Y=1047358
X732 169 175 177 3460 2 4 3477 ADDFHX1 $T=1385340 1027600 0 180 $X=1370160 $Y=1022160
X733 181 3506 176 3508 2 4 188 ADDFHX1 $T=1382040 1138480 1 0 $X=1382038 $Y=1133040
X734 3462 3558 3578 3582 2 4 3595 ADDFHX1 $T=1399860 1088080 0 0 $X=1399858 $Y=1087678
X735 162 3567 186 3579 2 4 3701 ADDFHX1 $T=1415040 1037680 0 0 $X=1415038 $Y=1037278
X736 5743 5730 5715 5592 2 4 5689 ADDFHX1 $T=2066460 1118320 0 180 $X=2051280 $Y=1112880
X737 5745 5732 5716 5648 2 4 5714 ADDFHX1 $T=2067120 1088080 0 180 $X=2051940 $Y=1082640
X738 385 6029 6007 6005 2 4 6001 ADDFHX1 $T=2160840 1047760 1 180 $X=2145660 $Y=1047358
X739 396 6135 6086 6110 2 4 6113 ADDFHX1 $T=2200440 1088080 1 180 $X=2185260 $Y=1087678
X740 402 6203 6192 399 2 4 6185 ADDFHX1 $T=2220900 1007440 0 180 $X=2205720 $Y=1002000
X741 2543 4 2548 2 2551 2560 NAND3X1 $T=1078440 1128400 1 0 $X=1078438 $Y=1122960
X742 3196 4 3212 2 3213 3178 NAND3X1 $T=1278420 1017520 0 0 $X=1278418 $Y=1017118
X743 4436 4 239 2 4420 238 NAND3X1 $T=1673760 1017520 1 0 $X=1673758 $Y=1012080
X744 6350 4 6339 2 6338 6247 NAND3X1 $T=2263140 1057840 0 180 $X=2260500 $Y=1052400
X745 5642 5628 5608 4 5578 2 AOI2BB1X2 $T=2036100 1088080 1 180 $X=2031480 $Y=1087678
X746 3477 3505 3523 3526 2 4 3531 ADDFHX2 $T=1376100 1007440 0 0 $X=1376098 $Y=1007038
X747 176 3515 3527 3528 2 4 3594 ADDFHX2 $T=1377420 1037680 1 0 $X=1377418 $Y=1032240
X748 3500 170 175 3519 2 4 3506 ADDFHX2 $T=1382700 1118320 1 0 $X=1382698 $Y=1112880
X749 3520 3453 162 3580 2 4 3593 ADDFHX2 $T=1393920 1057840 0 0 $X=1393918 $Y=1057438
X750 186 3528 190 3622 2 4 3633 ADDFHX2 $T=1409760 1027600 1 0 $X=1409758 $Y=1022160
X751 3579 3531 3633 3635 2 4 3638 ADDFHX2 $T=1411740 1017520 1 0 $X=1411738 $Y=1012080
X752 3594 3580 3701 3704 2 4 3713 ADDFHX2 $T=1431540 1047760 0 0 $X=1431538 $Y=1047358
X753 358 354 352 5732 2 4 5760 ADDFHX2 $T=2091540 1088080 1 180 $X=2069100 $Y=1087678
X754 353 356 5760 5767 2 4 350 ADDFHX2 $T=2092200 1128400 0 180 $X=2069760 $Y=1122960
X755 359 355 353 5730 2 4 5716 ADDFHX2 $T=2092200 1138480 0 180 $X=2069760 $Y=1133040
X756 6026 6012 6001 6004 2 4 5891 ADDFHX2 $T=2167440 1017520 0 180 $X=2145000 $Y=1012080
X757 6002 6005 6057 6041 2 4 6009 ADDFHX2 $T=2145660 1057840 0 0 $X=2145658 $Y=1057438
X758 6110 6126 6184 6149 2 4 6040 ADDFHX2 $T=2183280 1027600 1 0 $X=2183278 $Y=1022160
X759 4038 3317 4 2 4101 OR2X1 $T=1570800 1007440 1 0 $X=1570798 $Y=1002000
X760 119 2 88 4 CLKINVX3 $T=1144440 1108240 0 180 $X=1142460 $Y=1102800
X761 3259 2 3317 4 CLKINVX3 $T=1308120 1007440 1 0 $X=1308118 $Y=1002000
X762 3318 2 3366 4 CLKINVX3 $T=1333200 1027600 0 0 $X=1333198 $Y=1027198
X763 3825 2 3839 4 CLKINVX3 $T=1495560 1047760 1 0 $X=1495558 $Y=1042320
X764 4052 2 4037 4 CLKINVX3 $T=1558260 1078000 0 0 $X=1558258 $Y=1077598
X765 268 2 4852 4 CLKINVX3 $T=1792560 1118320 0 0 $X=1792558 $Y=1117918
X766 4855 2 4817 4 CLKINVX3 $T=1804440 1047760 1 0 $X=1804438 $Y=1042320
X767 5492 2 5482 4 CLKINVX3 $T=1991880 997360 1 180 $X=1989900 $Y=996958
X768 5503 2 4782 4 CLKINVX3 $T=1997160 1007440 0 180 $X=1995180 $Y=1002000
X769 403 2 410 4 CLKINVX3 $T=2230800 1088080 0 0 $X=2230798 $Y=1087678
X770 2281 2278 2 4 2259 AND2X1 $T=993300 1098160 1 180 $X=990660 $Y=1097758
X771 2175 2268 2 4 2323 AND2X1 $T=995940 1057840 1 0 $X=995938 $Y=1052400
X772 98 99 2 4 2576 AND2X1 $T=1104180 1007440 0 180 $X=1101540 $Y=1002000
X773 120 119 2 4 2556 AND2X1 $T=1146420 1078000 0 180 $X=1143780 $Y=1072560
X774 3141 3211 2 4 3297 AND2X1 $T=1298880 1037680 1 0 $X=1298878 $Y=1032240
X775 3209 3245 2 4 3273 AND2X1 $T=1301520 1078000 1 0 $X=1301518 $Y=1072560
X776 219 4311 2 4 220 AND2X1 $T=1636800 1057840 0 180 $X=1634160 $Y=1052400
X777 227 4311 2 4 223 AND2X1 $T=1642080 1007440 0 180 $X=1639440 $Y=1002000
X778 5410 5424 2 4 5441 AND2X1 $T=1976700 1118320 1 180 $X=1974060 $Y=1117918
X779 5668 5681 5664 2 5612 4 AOI2BB1X4 $T=2046660 1027600 1 180 $X=2039400 $Y=1027198
X780 283 280 2 284 4992 4922 4 AOI22X1 $T=1836120 1037680 1 0 $X=1836118 $Y=1032240
X781 283 281 2 284 4977 4964 4 AOI22X1 $T=1839420 1057840 1 180 $X=1836120 $Y=1057438
X782 283 279 2 284 5002 4976 4 AOI22X1 $T=1838760 1047760 0 0 $X=1838758 $Y=1047358
X783 283 295 2 284 5016 5118 4 AOI22X1 $T=1877700 1037680 0 180 $X=1874400 $Y=1032240
X784 313 283 2 5264 284 5172 4 AOI22X1 $T=1917960 1037680 0 180 $X=1914660 $Y=1032240
X785 315 283 2 312 284 5244 4 AOI22X1 $T=1917960 1037680 1 180 $X=1914660 $Y=1037278
X786 283 318 2 284 5162 5286 4 AOI22X1 $T=1925880 1037680 0 180 $X=1922580 $Y=1032240
X787 283 324 2 284 5274 5328 4 AOI22X1 $T=1944360 1037680 0 180 $X=1941060 $Y=1032240
X788 420 6583 2 6452 6363 6564 4 AOI22X1 $T=2352240 1128400 1 180 $X=2348940 $Y=1127998
X789 6675 6687 2 6486 6525 6676 4 AOI22X1 $T=2393820 1098160 0 180 $X=2390520 $Y=1092720
X790 389 407 353 6261 4 2 6263 ADDFXL $T=2226180 1047760 0 0 $X=2226178 $Y=1047358
X791 51 55 4 2 2004 XNOR2XL $T=921360 987280 0 180 $X=916080 $Y=981840
X792 3264 3292 4 2 3305 XNOR2XL $T=1301520 1088080 0 0 $X=1301518 $Y=1087678
X793 3713 3604 3714 2 4 OR2X4 $T=1456620 1067920 1 0 $X=1456618 $Y=1062480
X794 3908 3463 3920 2 4 OR2X4 $T=1519320 1047760 0 0 $X=1519318 $Y=1047358
X795 3909 3451 3942 2 4 OR2X4 $T=1525920 1088080 0 0 $X=1525918 $Y=1087678
X796 1901 4118 4128 2 4 OR2X4 $T=1579380 1078000 1 0 $X=1579378 $Y=1072560
X797 4326 4384 4388 2 4 OR2X4 $T=1655940 1088080 1 0 $X=1655938 $Y=1082640
X798 4267 4782 4801 2 4 OR2X4 $T=1776060 1017520 0 0 $X=1776058 $Y=1017118
X799 299 304 5142 2 4 OR2X4 $T=1887600 1138480 1 0 $X=1887598 $Y=1133040
X800 335 334 5457 2 4 OR2X4 $T=1994520 1138480 0 180 $X=1990560 $Y=1133040
X801 451 7149 7049 2 4 OR2X4 $T=2546280 1128400 0 180 $X=2542320 $Y=1122960
X802 63 67 4 2 INVX8 $T=978120 1118320 0 180 $X=974160 $Y=1112880
X803 5880 369 4 2 INVX8 $T=2112000 987280 0 180 $X=2108040 $Y=981840
X804 6041 6040 377 4 382 381 2 OAI2BB2X4 $T=2162160 987280 1 180 $X=2152260 $Y=986878
X805 1775 1805 1821 4 2 NAND2BX2 $T=850080 1078000 0 0 $X=850078 $Y=1077598
X806 4190 4170 4234 4 2 NAND2BX2 $T=1609740 1118320 1 180 $X=1605780 $Y=1117918
X807 4221 4128 4239 4 2 NAND2BX2 $T=1607100 1078000 0 0 $X=1607098 $Y=1077598
X808 47 2018 2017 1916 2 4 OAI2BB1X2 $T=909480 1088080 1 180 $X=904860 $Y=1087678
X809 3167 3091 3154 3166 2 4 OAI2BB1X2 $T=1264560 1007440 0 180 $X=1259940 $Y=1002000
X810 1795 1790 1849 4 2 NOR2BX2 $T=841500 1067920 0 0 $X=841498 $Y=1067518
X811 1792 1769 41 4 2 NOR2BX2 $T=842160 1128400 1 0 $X=842158 $Y=1122960
X812 4130 4106 4151 4 2 NOR2BX2 $T=1582020 1108240 0 0 $X=1582018 $Y=1107838
X813 3242 3297 4 2 3318 XOR2XL $T=1304160 1037680 1 0 $X=1304158 $Y=1032240
X814 4434 4547 4 2 4512 XOR2XL $T=1704780 1027600 0 180 $X=1699500 $Y=1022160
X815 236 235 4434 4442 232 2 4 219 SDFFRHQXL $T=1680360 1027600 1 180 $X=1663860 $Y=1027198
X816 236 235 4607 4600 232 2 4 4434 SDFFRHQXL $T=1729200 1037680 0 180 $X=1712700 $Y=1032240
X817 236 235 245 4592 232 2 4 250 SDFFRHQXL $T=1713360 1007440 1 0 $X=1713358 $Y=1002000
X818 236 277 279 4978 290 2 4 4977 SDFFRHQXL $T=1828860 1108240 0 0 $X=1828858 $Y=1107838
X819 236 277 280 4980 290 2 4 5008 SDFFRHQXL $T=1829520 1037680 0 0 $X=1829518 $Y=1037278
X820 236 277 4977 4981 290 2 4 5002 SDFFRHQXL $T=1829520 1078000 0 0 $X=1829518 $Y=1077598
X821 236 277 250 4982 290 2 4 5021 SDFFRHQXL $T=1832160 1007440 0 0 $X=1832158 $Y=1007038
X822 236 277 281 4923 290 2 4 5019 SDFFRHQXL $T=1832160 1017520 0 0 $X=1832158 $Y=1017118
X823 236 277 4992 5082 290 2 4 5016 SDFFRHQXL $T=1867800 1037680 1 180 $X=1851300 $Y=1037278
X824 236 277 5002 5066 290 2 4 4992 SDFFRHQXL $T=1855260 1057840 0 0 $X=1855258 $Y=1057438
X825 236 277 5016 5083 290 2 4 5132 SDFFRHQXL $T=1859880 1017520 1 0 $X=1859878 $Y=1012080
X826 236 277 295 5203 290 2 4 5162 SDFFRHQXL $T=1902780 1017520 1 180 $X=1886280 $Y=1017118
X827 236 277 5162 5182 290 2 4 5238 SDFFRHQXL $T=1886940 1007440 0 0 $X=1886938 $Y=1007038
X828 236 277 5274 5295 290 2 4 5264 SDFFRHQXL $T=1928520 1047760 1 180 $X=1912020 $Y=1047358
X829 236 277 313 5245 290 2 4 5326 SDFFRHQXL $T=1914000 1017520 1 0 $X=1913998 $Y=1012080
X830 236 277 5264 320 290 2 4 5384 SDFFRHQXL $T=1934460 1088080 1 0 $X=1934458 $Y=1082640
X831 236 277 324 5367 290 2 4 5274 SDFFRHQXL $T=1954260 1047760 1 180 $X=1937760 $Y=1047358
X832 236 277 318 5323 290 2 4 5387 SDFFRHQXL $T=1938420 1017520 0 0 $X=1938418 $Y=1017118
X833 236 277 315 5354 290 2 4 5398 SDFFRHQXL $T=1940400 1017520 1 0 $X=1940398 $Y=1012080
X834 5021 2 281 4 BUFX3 $T=1841400 1007440 0 180 $X=1838760 $Y=1002000
X835 5019 2 280 4 BUFX3 $T=1841400 1027600 0 180 $X=1838760 $Y=1022160
X836 5008 2 279 4 BUFX3 $T=1845360 1037680 0 180 $X=1842720 $Y=1032240
X837 5132 2 295 4 BUFX3 $T=1875720 1007440 0 180 $X=1873080 $Y=1002000
X838 316 2 311 4 BUFX3 $T=1915980 1118320 1 180 $X=1913340 $Y=1117918
X839 5238 2 313 4 BUFX3 $T=1914660 1007440 0 0 $X=1914658 $Y=1007038
X840 5326 2 315 4 BUFX3 $T=1933140 997360 0 0 $X=1933138 $Y=996958
X841 5398 2 318 4 BUFX3 $T=1954260 1007440 0 180 $X=1951620 $Y=1002000
X842 5384 2 332 4 BUFX3 $T=1959540 1088080 1 0 $X=1959538 $Y=1082640
X843 5387 2 324 4 BUFX3 $T=1962180 1017520 0 0 $X=1962178 $Y=1017118
X844 347 2 383 4 BUFX3 $T=2245980 1138480 1 0 $X=2245978 $Y=1133040
X845 3015 2796 4 2 3017 3058 AOI2BB1X1 $T=1225620 997360 0 0 $X=1225618 $Y=996958
X846 282 4991 2 285 287 4977 4974 288 4 AOI222X1 $T=1836780 1128400 1 0 $X=1836778 $Y=1122960
X847 4993 282 2 286 287 5002 4994 288 4 AOI222X1 $T=1837440 1098160 0 0 $X=1837438 $Y=1097758
X848 5087 282 2 5065 287 4992 5064 288 4 AOI222X1 $T=1859880 1078000 0 180 $X=1854600 $Y=1072560
X849 5151 282 2 5152 287 5016 5141 288 4 AOI222X1 $T=1883640 1067920 1 180 $X=1878360 $Y=1067518
X850 5234 282 2 5202 287 5162 5195 288 4 AOI222X1 $T=1900800 1067920 1 180 $X=1895520 $Y=1067518
X851 5279 282 2 5324 287 288 5327 5264 4 AOI222X1 $T=1933140 1067920 1 180 $X=1927860 $Y=1067518
X852 5278 282 2 5337 287 5274 5336 288 4 AOI222X1 $T=1942380 1067920 1 180 $X=1937100 $Y=1067518
X853 123 2786 2795 4 2 127 XNOR3X2 $T=1155000 997360 1 0 $X=1154998 $Y=991920
X854 3015 2885 2796 4 2 3091 XNOR3X2 $T=1231560 1007440 1 0 $X=1231558 $Y=1002000
X855 155 3118 3105 4 2 3226 XNOR3X2 $T=1251360 1118320 0 0 $X=1251358 $Y=1117918
X856 3154 3241 3091 4 2 3259 XNOR3X2 $T=1281720 1007440 0 0 $X=1281718 $Y=1007038
X857 233 2 234 230 228 4405 4 AOI22XL $T=1661220 997360 1 0 $X=1661218 $Y=991920
X858 233 2 4403 230 219 4406 4 AOI22XL $T=1661220 1047760 1 0 $X=1661218 $Y=1042320
X859 233 2 4512 230 4434 4564 4 AOI22XL $T=1700160 1037680 1 0 $X=1700158 $Y=1032240
X860 233 2 4544 230 245 4577 4 AOI22XL $T=1710720 987280 0 0 $X=1710718 $Y=986878
X861 233 2 4545 230 250 4575 4 AOI22XL $T=1712700 1017520 0 0 $X=1712698 $Y=1017118
X862 374 398 4 2 BUFX4 $T=2259180 1098160 0 0 $X=2259178 $Y=1097758
X863 4578 4576 4 2 4548 NAND2BX4 $T=1715340 1067920 0 180 $X=1710060 $Y=1062480
X864 219 4309 221 2 4 222 OR3XL $T=1634160 987280 1 0 $X=1634158 $Y=981840
X865 228 227 229 2 4 4309 OR3XL $T=1657920 987280 1 180 $X=1654620 $Y=986878
X866 46 48 49 4 50 2 2003 OAI31X1 $T=899580 987280 1 0 $X=899578 $Y=981840
X867 3166 3178 3176 3194 4 2 AND3X4 $T=1268520 1007440 1 0 $X=1268518 $Y=1002000
X868 2 219 224 225 4309 226 4 NOR4X1 $T=1640100 987280 0 0 $X=1640098 $Y=986878
X869 2 222 242 244 247 4436 4 NOR4X1 $T=1681680 987280 1 0 $X=1681678 $Y=981840
X870 2 4977 5002 4992 5016 5051 4 NOR4X1 $T=1844040 1057840 0 0 $X=1844038 $Y=1057438
X871 2 4977 5002 4992 5016 5006 4 NOR4X1 $T=1844040 1067920 1 0 $X=1844038 $Y=1062480
X872 2 5162 5274 5264 312 5007 4 NOR4X1 $T=1918620 1057840 1 180 $X=1914660 $Y=1057438
X873 2 5162 5274 5264 312 5267 4 NOR4X1 $T=1922580 1057840 0 0 $X=1922578 $Y=1057438
X874 4434 4 4420 2 4436 237 NAND3XL $T=1670460 1017520 0 180 $X=1667820 $Y=1012080
X875 4436 4 239 2 245 243 NAND3XL $T=1682340 1017520 1 0 $X=1682338 $Y=1012080
X876 300 4 296 2 274 5131 NAND3XL $T=1878360 987280 0 180 $X=1875720 $Y=981840
X877 300 296 301 4 5138 2 OAI2BB1XL $T=1886940 987280 0 180 $X=1883640 $Y=981840
X878 3194 4 157 2 CLKINVX8 $T=1272480 1007440 1 0 $X=1272478 $Y=1002000
X879 236 235 260 4589 232 4607 4 2 261 SDFFRXL $T=1711380 1098160 1 0 $X=1711378 $Y=1092720
X880 236 235 264 4621 232 260 4 2 262 SDFFRXL $T=1723260 1118320 0 0 $X=1723258 $Y=1117918
X881 6969 4384 4 2 BUFX16 $T=2498760 1098160 1 0 $X=2498758 $Y=1092720
X882 236 235 219 4410 232 2 4 228 SDFFRHQX1 $T=1669800 1007440 0 180 $X=1653300 $Y=1002000
X883 236 235 248 4606 232 2 4 245 SDFFRHQX1 $T=1729860 997360 1 180 $X=1713360 $Y=996958
X884 6934 4360 4 2 BUFX12 $T=2484240 1108240 0 0 $X=2484238 $Y=1107838
X885 444 4421 4 2 BUFX12 $T=2500080 1138480 1 0 $X=2500078 $Y=1133040
X886 251 4 250 248 245 246 2 NAND4X1 $T=1687620 997360 0 180 $X=1684320 $Y=991920
X887 3195 3209 4 3198 3197 3177 2 AOI2BB2X2 $T=1279740 1047760 1 180 $X=1273800 $Y=1047358
X888 229 228 224 225 4 2 4311 AND4X2 $T=1651320 987280 1 180 $X=1647360 $Y=986878
X889 3216 158 4 159 3226 160 3230 3213 2 OAI222X2 $T=1278420 1118320 1 0 $X=1278418 $Y=1112880
X890 3216 158 4 159 3226 161 3230 3264 2 OAI222X2 $T=1304160 1118320 1 0 $X=1304158 $Y=1112880
X891 4420 2 248 250 4434 252 4 NOR4BXL $T=1684320 997360 0 0 $X=1684318 $Y=996958
X892 400 358 401 6228 4 2 6215 ADDFX1 $T=2209680 1088080 1 0 $X=2209678 $Y=1082640
.ENDS
***************************************
.SUBCKT NAND4BBX1 BN D C VDD AN Y VSS
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3BX4 AN C VSS B Y VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR3XL C VDD B VSS A Y
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFSXL CK SE SI D SN QN VSS VDD Q
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX4 A Y VSS VDD
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4XL D VSS C B Y A VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI222XL C0 C1 VDD B1 B0 A0 A1 Y VSS
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX1 A VSS VDD Y
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB2X4 A0N A1N B0 VSS B1 Y VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR4X4 A B C D Y VSS VDD
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB2XL A0N A1N B1 B0 VSS VDD Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_61 1 3 5 7 22 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39
+ 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
+ 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79
+ 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99
+ 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119
+ 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139
+ 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159
+ 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179
+ 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199
+ 200 201 202 203 204 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 531 532 533 534 535 536 537 538 539 540 541 542 543
+ 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563
+ 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583
+ 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603
+ 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623
+ 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643
+ 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663
+ 664 665 666 667 668 669 670 671 672 673 675 676 677 678 679 680 681 682 684 685
+ 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 701 702 703 704 705
+ 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723 724 725
+ 726 727 728 729 730 731 732 733 734 735 736 737 738 739 740 741 742 743 744 745
+ 746 747 748 749 750 751 752 753 754 755 756 757 779 1548 1549
** N=26792 EP=735 IP=11689 FDC=0
X0 3996 200 3 1 BUFX20 $T=1283040 1561840 0 180 $X=1272480 $Y=1556400
X1 25 1 27 3 30 NAND2X1 $T=661320 1511440 1 0 $X=661318 $Y=1506000
X2 35 1 37 3 25 NAND2X1 $T=667920 1531600 0 0 $X=667918 $Y=1531198
X3 1598 1 1581 3 1593 NAND2X1 $T=675840 1541680 1 0 $X=675838 $Y=1536240
X4 53 1 1661 3 1654 NAND2X1 $T=693660 1541680 1 0 $X=693658 $Y=1536240
X5 59 1 1723 3 1721 NAND2X1 $T=704220 1582000 1 0 $X=704218 $Y=1576560
X6 1654 1 1735 3 1844 NAND2X1 $T=705540 1491280 0 0 $X=705538 $Y=1490878
X7 1721 1 1764 3 1780 NAND2X1 $T=716100 1491280 1 0 $X=716098 $Y=1485840
X8 1780 1 1565 3 1798 NAND2X1 $T=718740 1491280 1 0 $X=718738 $Y=1485840
X9 1805 1 1802 3 1742 NAND2X1 $T=726000 1602160 0 180 $X=724020 $Y=1596720
X10 1817 1 1850 3 1863 NAND2X1 $T=737220 1582000 1 0 $X=737218 $Y=1576560
X11 1878 1 1856 3 1814 NAND2X1 $T=745140 1461040 1 0 $X=745138 $Y=1455600
X12 1928 1 1930 3 1816 NAND2X1 $T=753720 1551760 0 0 $X=753718 $Y=1551358
X13 1997 1 1927 3 1862 NAND2X1 $T=760980 1450960 0 0 $X=760978 $Y=1450558
X14 1960 1 1959 3 1805 NAND2X1 $T=762300 1602160 1 0 $X=762298 $Y=1596720
X15 1993 1 1992 3 1875 NAND2X1 $T=770880 1551760 0 0 $X=770878 $Y=1551358
X16 2347 1 1961 3 2363 NAND2X1 $T=877140 1501360 0 180 $X=875160 $Y=1495920
X17 2363 1 2348 3 2379 NAND2X1 $T=878460 1511440 1 0 $X=878458 $Y=1506000
X18 2444 1 113 3 2479 NAND2X1 $T=898260 1602160 0 0 $X=898258 $Y=1601758
X19 1687 1 2476 3 2477 NAND2X1 $T=903540 1450960 1 0 $X=903538 $Y=1445520
X20 112 1 2479 3 2516 NAND2X1 $T=907500 1612240 0 0 $X=907498 $Y=1611838
X21 2500 1 1929 3 2515 NAND2X1 $T=910800 1481200 1 180 $X=908820 $Y=1480798
X22 2533 1 2534 3 2498 NAND2X1 $T=919380 1461040 1 180 $X=917400 $Y=1460638
X23 2707 1 2632 3 2621 NAND2X1 $T=948420 1471120 0 180 $X=946440 $Y=1465680
X24 125 1 126 3 2707 NAND2X1 $T=965580 1471120 1 180 $X=963600 $Y=1470718
X25 2834 1 2804 3 2805 NAND2X1 $T=982080 1602160 1 180 $X=980100 $Y=1601758
X26 2826 1 2772 3 2759 NAND2X1 $T=984720 1491280 1 180 $X=982740 $Y=1490878
X27 137 1 135 3 2826 NAND2X1 $T=993300 1481200 1 180 $X=991320 $Y=1480798
X28 140 1 141 3 2791 NAND2X1 $T=993300 1521520 1 0 $X=993298 $Y=1516080
X29 2904 1 2903 3 2832 NAND2X1 $T=1001220 1471120 0 0 $X=1001218 $Y=1470718
X30 147 1 150 3 151 NAND2X1 $T=1007820 1541680 1 0 $X=1007818 $Y=1536240
X31 154 1 152 3 2807 NAND2X1 $T=1011780 1602160 1 0 $X=1011778 $Y=1596720
X32 3142 1 3140 3 171 NAND2X1 $T=1067220 1481200 1 180 $X=1065240 $Y=1480798
X33 3158 1 177 3 3140 NAND2X1 $T=1069860 1481200 0 180 $X=1067880 $Y=1475760
X34 181 1 179 3 3127 NAND2X1 $T=1071180 1440880 0 180 $X=1069200 $Y=1435440
X35 3171 1 3159 3 3142 NAND2X1 $T=1075140 1481200 1 180 $X=1073160 $Y=1480798
X36 3190 1 3193 3 3177 NAND2X1 $T=1085040 1440880 0 0 $X=1085038 $Y=1440478
X37 3434 1 3390 3 3338 NAND2X1 $T=1133880 1511440 0 180 $X=1131900 $Y=1506000
X38 3408 1 3395 3 3356 NAND2X1 $T=1136520 1521520 1 180 $X=1134540 $Y=1521118
X39 3399 1 3397 3 3391 NAND2X1 $T=1137840 1461040 1 180 $X=1135860 $Y=1460638
X40 3429 1 3433 3 3520 NAND2X1 $T=1145100 1531600 1 0 $X=1145098 $Y=1526160
X41 3480 1 3492 3 3497 NAND2X1 $T=1155660 1501360 0 0 $X=1155658 $Y=1500958
X42 223 1 199 3 3553 NAND2X1 $T=1170840 1531600 1 0 $X=1170838 $Y=1526160
X43 3553 1 3556 3 3564 NAND2X1 $T=1172820 1531600 1 0 $X=1172818 $Y=1526160
X44 228 1 207 3 3556 NAND2X1 $T=1176120 1531600 1 0 $X=1176118 $Y=1526160
X45 3792 1 275 3 3837 NAND2X1 $T=1228260 1561840 1 0 $X=1228258 $Y=1556400
X46 279 1 3845 3 3840 NAND2X1 $T=1236840 1541680 0 0 $X=1236838 $Y=1541278
X47 290 1 3857 3 3882 NAND2X1 $T=1248060 1440880 1 0 $X=1248058 $Y=1435440
X48 293 1 3919 3 3924 NAND2X1 $T=1257300 1481200 0 0 $X=1257298 $Y=1480798
X49 3937 1 300 3 4134 NAND2X1 $T=1275780 1450960 0 0 $X=1275778 $Y=1450558
X50 305 1 3986 3 4017 NAND2X1 $T=1281060 1450960 1 0 $X=1281058 $Y=1445520
X51 328 1 3037 3 4057 NAND2X1 $T=1321320 1571920 0 180 $X=1319340 $Y=1566480
X52 85 1 4145 3 4143 NAND2X1 $T=1325280 1501360 1 180 $X=1323300 $Y=1500958
X53 345 1 2577 3 4394 NAND2X1 $T=1385340 1501360 0 180 $X=1383360 $Y=1495920
X54 4490 1 4488 3 4506 NAND2X1 $T=1409100 1571920 0 180 $X=1407120 $Y=1566480
X55 2518 1 350 3 4507 NAND2X1 $T=1409100 1521520 0 0 $X=1409098 $Y=1521118
X56 349 1 355 3 4530 NAND2X1 $T=1427580 1461040 0 0 $X=1427578 $Y=1460638
X57 4635 1 4577 3 4528 NAND2X1 $T=1434840 1450960 0 180 $X=1432860 $Y=1445520
X58 4487 1 4617 3 4581 NAND2X1 $T=1442100 1551760 0 0 $X=1442098 $Y=1551358
X59 4532 1 4637 3 4685 NAND2X1 $T=1453980 1511440 0 0 $X=1453978 $Y=1511038
X60 4704 1 4692 3 4691 NAND2X1 $T=1455960 1450960 0 180 $X=1453980 $Y=1445520
X61 4802 1 4727 3 4792 NAND2X1 $T=1479060 1531600 0 180 $X=1477080 $Y=1526160
X62 4583 1 4785 3 4726 NAND2X1 $T=1479060 1501360 1 0 $X=1479058 $Y=1495920
X63 376 1 4870 3 4854 NAND2X1 $T=1500840 1450960 1 0 $X=1500838 $Y=1445520
X64 4851 1 4779 3 4897 NAND2X1 $T=1500840 1541680 1 0 $X=1500838 $Y=1536240
X65 5022 1 5001 3 4227 NAND2X1 $T=1534500 1531600 0 180 $X=1532520 $Y=1526160
X66 5025 1 5001 3 4041 NAND2X1 $T=1541760 1531600 0 180 $X=1539780 $Y=1526160
X67 412 1 5240 3 5207 NAND2X1 $T=1584660 1592080 0 0 $X=1584658 $Y=1591678
X68 5247 1 5237 3 5239 NAND2X1 $T=1586640 1571920 0 180 $X=1584660 $Y=1566480
X69 5180 1 5357 3 419 NAND2X1 $T=1615680 1511440 1 0 $X=1615678 $Y=1506000
X70 5115 1 396 3 5112 NAND2X1 $T=1620960 1511440 1 0 $X=1620958 $Y=1506000
X71 411 1 5460 3 5461 NAND2X1 $T=1648020 1450960 1 180 $X=1646040 $Y=1450558
X72 5498 1 438 3 411 NAND2X1 $T=1650660 1501360 1 180 $X=1648680 $Y=1500958
X73 6159 1 6156 3 6139 NAND2X1 $T=1822260 1450960 0 180 $X=1820280 $Y=1445520
X74 6357 1 6288 3 6330 NAND2X1 $T=1870440 1602160 0 180 $X=1868460 $Y=1596720
X75 6494 1 6173 3 6442 NAND2X1 $T=1908060 1592080 1 180 $X=1906080 $Y=1591678
X76 6996 1 604 3 7050 NAND2X1 $T=2061840 1531600 1 0 $X=2061838 $Y=1526160
X77 7075 1 609 3 7069 NAND2X1 $T=2065140 1551760 1 180 $X=2063160 $Y=1551358
X78 557 1 567 3 7100 NAND2X1 $T=2075700 1511440 0 180 $X=2073720 $Y=1506000
X79 7120 1 7119 3 7108 NAND2X1 $T=2080980 1521520 0 180 $X=2079000 $Y=1516080
X80 568 1 7139 3 7132 NAND2X1 $T=2085600 1461040 1 0 $X=2085598 $Y=1455600
X81 623 1 624 3 7171 NAND2X1 $T=2124540 1582000 0 0 $X=2124538 $Y=1581598
X82 629 1 7342 3 7310 NAND2X1 $T=2141700 1531600 1 0 $X=2141698 $Y=1526160
X83 631 1 633 3 7328 NAND2X1 $T=2144340 1612240 1 0 $X=2144338 $Y=1606800
X84 636 1 635 3 7473 NAND2X1 $T=2153580 1440880 0 180 $X=2151600 $Y=1435440
X85 7442 1 7426 3 7427 NAND2X1 $T=2156880 1531600 0 180 $X=2154900 $Y=1526160
X86 638 1 7444 3 637 NAND2X1 $T=2158200 1602160 1 180 $X=2156220 $Y=1601758
X87 7443 1 7445 3 7429 NAND2X1 $T=2156880 1561840 0 0 $X=2156878 $Y=1561438
X88 639 1 7423 3 7368 NAND2X1 $T=2159520 1521520 1 180 $X=2157540 $Y=1521118
X89 7571 1 7528 3 7448 NAND2X1 $T=2179980 1461040 1 180 $X=2178000 $Y=1460638
X90 7548 1 7531 3 7488 NAND2X1 $T=2181300 1582000 0 180 $X=2179320 $Y=1576560
X91 7530 1 7490 3 7512 NAND2X1 $T=2183280 1561840 1 0 $X=2183278 $Y=1556400
X92 7557 1 7555 3 7442 NAND2X1 $T=2187900 1531600 0 180 $X=2185920 $Y=1526160
X93 7467 1 7528 3 7570 NAND2X1 $T=2199120 1471120 0 0 $X=2199118 $Y=1470718
X94 7649 1 647 3 7571 NAND2X1 $T=2201100 1461040 0 180 $X=2199120 $Y=1455600
X95 7670 1 648 3 7397 NAND2X1 $T=2209020 1461040 1 0 $X=2209018 $Y=1455600
X96 650 1 7712 3 7648 NAND2X1 $T=2216280 1521520 1 0 $X=2216278 $Y=1516080
X97 7727 1 7729 3 7693 NAND2X1 $T=2225520 1592080 1 0 $X=2225518 $Y=1586640
X98 7772 1 7757 3 7726 NAND2X1 $T=2234100 1571920 1 180 $X=2232120 $Y=1571518
X99 7788 1 655 3 7766 NAND2X1 $T=2238720 1450960 0 180 $X=2236740 $Y=1445520
X100 654 1 7791 3 7772 NAND2X1 $T=2238060 1592080 0 0 $X=2238058 $Y=1591678
X101 7757 1 7815 3 7804 NAND2X1 $T=2245320 1582000 0 0 $X=2245318 $Y=1581598
X102 660 1 7881 3 7880 NAND2X1 $T=2261820 1582000 0 0 $X=2261818 $Y=1581598
X103 7913 1 662 3 7894 NAND2X1 $T=2266440 1461040 0 180 $X=2264460 $Y=1455600
X104 7945 1 7946 3 7882 NAND2X1 $T=2280300 1531600 1 0 $X=2280298 $Y=1526160
X105 7972 1 7862 3 7899 NAND2X1 $T=2285580 1531600 0 0 $X=2285578 $Y=1531198
X106 7974 1 7980 3 7972 NAND2X1 $T=2292180 1541680 0 0 $X=2292178 $Y=1541278
X107 675 1 672 3 7958 NAND2X1 $T=2303400 1612240 1 180 $X=2301420 $Y=1611838
X108 673 1 7990 3 8068 NAND2X1 $T=2309340 1571920 0 0 $X=2309338 $Y=1571518
X109 8089 1 8062 3 8087 NAND2X1 $T=2313960 1511440 0 180 $X=2311980 $Y=1506000
X110 8119 1 8101 3 8089 NAND2X1 $T=2322540 1521520 0 0 $X=2322538 $Y=1521118
X111 8137 1 8200 3 8208 NAND2X1 $T=2348280 1521520 1 0 $X=2348278 $Y=1516080
X112 8247 1 8245 3 8199 NAND2X1 $T=2359500 1521520 1 180 $X=2357520 $Y=1521118
X113 8244 1 694 3 8186 NAND2X1 $T=2364120 1440880 1 0 $X=2364118 $Y=1435440
X114 8345 1 8353 3 8347 NAND2X1 $T=2403060 1481200 0 0 $X=2403058 $Y=1480798
X115 8511 1 8508 3 8478 NAND2X1 $T=2428800 1481200 1 180 $X=2426820 $Y=1480798
X116 8560 1 8424 3 708 NAND2X1 $T=2442000 1440880 0 180 $X=2440020 $Y=1435440
X117 8627 1 8551 3 8558 NAND2X1 $T=2458500 1481200 1 0 $X=2458498 $Y=1475760
X118 8671 1 8682 3 714 NAND2X1 $T=2478960 1461040 0 0 $X=2478958 $Y=1460638
X119 8786 1 718 3 716 NAND2X1 $T=2488860 1430800 1 180 $X=2486880 $Y=1430398
X120 8883 1 8781 3 731 NAND2X1 $T=2523840 1450960 1 0 $X=2523838 $Y=1445520
X121 8884 1 8910 3 8882 NAND2X1 $T=2536380 1450960 1 0 $X=2536378 $Y=1445520
X122 9046 1 9084 3 741 NAND2X1 $T=2572020 1430800 1 180 $X=2570040 $Y=1430398
X123 9117 1 742 3 745 NAND2X1 $T=2578620 1440880 0 0 $X=2578618 $Y=1440478
X124 9220 1 9236 3 752 NAND2X1 $T=2605680 1450960 1 0 $X=2605678 $Y=1445520
X125 2421 3 1 111 2395 NOR2X4 $T=894960 1531600 0 180 $X=890340 $Y=1526160
X126 134 3 1 131 2723 NOR2X4 $T=985380 1440880 0 0 $X=985378 $Y=1440478
X127 3564 3 1 3588 238 NOR2X4 $T=1181400 1531600 1 0 $X=1181398 $Y=1526160
X128 313 3 1 3883 4054 NOR2X4 $T=1301520 1531600 1 180 $X=1296900 $Y=1531198
X129 4097 3 1 4086 3996 NOR2X4 $T=1310100 1561840 0 180 $X=1305480 $Y=1556400
X130 336 3 1 2604 4305 NOR2X4 $T=1361580 1561840 0 180 $X=1356960 $Y=1556400
X131 4728 3 1 4723 4729 NOR2X4 $T=1463880 1602160 0 180 $X=1459260 $Y=1596720
X132 4729 3 1 4753 4780 NOR2X4 $T=1466520 1602160 0 0 $X=1466518 $Y=1601758
X133 4744 3 1 4745 4753 NOR2X4 $T=1475100 1612240 0 180 $X=1470480 $Y=1606800
X134 4510 3 1 4855 4800 NOR2X4 $T=1498200 1481200 0 0 $X=1498198 $Y=1480798
X135 5151 3 1 4831 5176 NOR2X4 $T=1568820 1592080 1 180 $X=1564200 $Y=1591678
X136 5696 3 1 5625 5626 NOR2X4 $T=1707420 1491280 0 180 $X=1702800 $Y=1485840
X137 5748 3 1 5255 5726 NOR2X4 $T=1721280 1491280 1 180 $X=1716660 $Y=1490878
X138 5496 3 1 5255 5698 NOR2X4 $T=1725240 1491280 0 0 $X=1725238 $Y=1490878
X139 6705 3 1 580 6721 NOR2X4 $T=1970760 1531600 0 180 $X=1966140 $Y=1526160
X140 581 3 1 578 6666 NOR2X4 $T=1968780 1521520 1 0 $X=1968778 $Y=1516080
X141 6756 3 1 6787 6818 NOR2X4 $T=1987920 1481200 1 0 $X=1987918 $Y=1475760
X142 6779 3 1 590 6787 NOR2X4 $T=1989900 1501360 0 0 $X=1989898 $Y=1500958
X143 601 3 1 6944 6946 NOR2X4 $T=2034120 1491280 0 0 $X=2034118 $Y=1490878
X144 6974 3 1 600 6930 NOR2X4 $T=2036100 1511440 1 0 $X=2036098 $Y=1506000
X145 7372 3 1 7306 7360 NOR2X4 $T=2146320 1511440 1 180 $X=2141700 $Y=1511038
X146 639 3 1 7423 7365 NOR2X4 $T=2157540 1511440 0 0 $X=2157538 $Y=1511038
X147 663 3 1 7926 7794 NOR2X4 $T=2269740 1491280 0 0 $X=2269738 $Y=1490878
X148 7 1 26 1605 3 NAND2BX1 $T=661320 1450960 0 0 $X=661318 $Y=1450558
X149 1818 1 1814 1738 3 NAND2BX1 $T=730620 1461040 0 180 $X=727980 $Y=1455600
X150 1819 1 1816 1767 3 NAND2BX1 $T=730620 1561840 0 180 $X=727980 $Y=1556400
X151 2723 1 2725 2700 3 NAND2BX1 $T=962940 1440880 1 180 $X=960300 $Y=1440478
X152 2781 1 2791 2624 3 NAND2BX1 $T=982740 1521520 1 180 $X=980100 $Y=1521118
X153 2819 1 2807 2806 3 NAND2BX1 $T=982740 1602160 0 180 $X=980100 $Y=1596720
X154 2837 1 138 2804 3 NAND2BX1 $T=990660 1612240 0 180 $X=988020 $Y=1606800
X155 2837 1 2834 132 3 NAND2BX1 $T=990660 1612240 1 180 $X=988020 $Y=1611838
X156 2973 1 2970 2907 3 NAND2BX1 $T=1023000 1491280 0 180 $X=1020360 $Y=1485840
X157 312 1 311 4040 3 NAND2BX1 $T=1298220 1491280 1 180 $X=1295580 $Y=1490878
X158 312 1 311 4036 3 NAND2BX1 $T=1298880 1501360 0 180 $X=1296240 $Y=1495920
X159 4305 1 4289 4351 3 NAND2BX1 $T=1366860 1551760 1 0 $X=1366858 $Y=1546320
X160 4368 1 4353 4404 3 NAND2BX1 $T=1377420 1561840 0 0 $X=1377418 $Y=1561438
X161 4522 1 4506 4544 3 NAND2BX1 $T=1418340 1561840 0 0 $X=1418338 $Y=1561438
X162 4560 1 4581 4508 3 NAND2BX1 $T=1435500 1551760 1 180 $X=1432860 $Y=1551358
X163 4784 1 4726 4720 3 NAND2BX1 $T=1463880 1491280 1 180 $X=1461240 $Y=1490878
X164 4800 1 4815 4801 3 NAND2BX1 $T=1490280 1471120 0 180 $X=1487640 $Y=1465680
X165 5496 1 466 5748 3 NAND2BX1 $T=1721280 1491280 0 180 $X=1718640 $Y=1485840
X166 567 1 568 6600 3 NAND2BX1 $T=1939740 1511440 0 0 $X=1939738 $Y=1511038
X167 614 1 613 7131 3 NAND2BX1 $T=2086260 1440880 0 180 $X=2083620 $Y=1435440
X168 7365 1 7368 7290 3 NAND2BX1 $T=2151600 1521520 0 180 $X=2148960 $Y=1516080
X169 641 1 7473 7549 3 NAND2BX1 $T=2180640 1430800 0 0 $X=2180638 $Y=1430398
X170 7531 1 644 7443 3 NAND2BX1 $T=2183280 1571920 0 0 $X=2183278 $Y=1571518
X171 7668 1 7648 7529 3 NAND2BX1 $T=2203080 1511440 1 180 $X=2200440 $Y=1511038
X172 7711 1 7707 7650 3 NAND2BX1 $T=2216940 1501360 0 180 $X=2214300 $Y=1495920
X173 649 1 7757 7684 3 NAND2BX1 $T=2231460 1592080 1 180 $X=2228820 $Y=1591678
X174 7783 1 7766 7756 3 NAND2BX1 $T=2232780 1450960 1 180 $X=2230140 $Y=1450558
X175 7893 1 7894 7875 3 NAND2BX1 $T=2264460 1471120 0 180 $X=2261820 $Y=1465680
X176 7794 1 7864 7751 3 NAND2BX1 $T=2267100 1491280 0 180 $X=2264460 $Y=1485840
X177 669 1 672 7997 3 NAND2BX1 $T=2291520 1612240 1 0 $X=2291518 $Y=1606800
X178 8144 1 8121 8053 3 NAND2BX1 $T=2325840 1511440 1 180 $X=2323200 $Y=1511038
X179 8228 1 8199 8167 3 NAND2BX1 $T=2350260 1491280 0 180 $X=2347620 $Y=1485840
X180 8265 1 8275 8262 3 NAND2BX1 $T=2374020 1511440 1 0 $X=2374018 $Y=1506000
X181 8351 1 8347 8292 3 NAND2BX1 $T=2389860 1461040 0 180 $X=2387220 $Y=1455600
X182 8421 1 8428 8357 3 NAND2BX1 $T=2404380 1471120 1 180 $X=2401740 $Y=1470718
X183 8561 1 8558 707 3 NAND2BX1 $T=2445960 1461040 1 180 $X=2443320 $Y=1460638
X184 63 1840 1 1805 3 1823 OAI21X1 $T=739860 1602160 1 0 $X=739858 $Y=1596720
X185 1814 1872 1 1862 3 71 OAI21X1 $T=744480 1450960 1 0 $X=744478 $Y=1445520
X186 2724 2781 1 2791 3 2762 OAI21X1 $T=975480 1521520 1 0 $X=975478 $Y=1516080
X187 2834 2819 1 2807 3 2827 OAI21X1 $T=997260 1602160 0 180 $X=993960 $Y=1596720
X188 2918 2938 1 2948 3 158 OAI21X1 $T=1019700 1481200 0 180 $X=1016400 $Y=1475760
X189 157 156 1 160 3 2954 OAI21X1 $T=1017720 1440880 0 0 $X=1017718 $Y=1440478
X190 4353 4305 1 4289 3 4347 OAI21X1 $T=1373460 1551760 1 180 $X=1370160 $Y=1551358
X191 4868 4856 1 328 3 4688 OAI21X1 $T=1498860 1571920 0 180 $X=1495560 $Y=1566480
X192 4897 359 1 4898 3 380 OAI21X1 $T=1500840 1531600 1 0 $X=1500838 $Y=1526160
X193 7331 7312 1 7310 3 7289 OAI21X1 $T=2132460 1521520 1 180 $X=2129160 $Y=1521118
X194 7365 7310 1 7368 3 7372 OAI21X1 $T=2142360 1521520 1 0 $X=2142358 $Y=1516080
X195 641 642 1 7473 3 7472 OAI21X1 $T=2169420 1430800 1 180 $X=2166120 $Y=1430398
X196 7711 7608 1 7707 3 7748 OAI21X1 $T=2223540 1491280 0 0 $X=2223538 $Y=1490878
X197 43 1 25 1593 3 46 OAI21XL $T=673860 1521520 0 0 $X=673858 $Y=1521118
X198 1760 1 44 1659 3 1739 OAI21XL $T=710820 1511440 1 180 $X=708180 $Y=1511038
X199 1819 1 1765 1816 3 1813 OAI21XL $T=729960 1551760 1 180 $X=727320 $Y=1551358
X200 1848 1 44 1834 3 68 OAI21XL $T=733920 1511440 1 180 $X=731280 $Y=1511038
X201 1822 1 44 1782 3 1945 OAI21XL $T=739200 1511440 1 0 $X=739198 $Y=1506000
X202 1816 1 1849 1875 3 1826 OAI21XL $T=743160 1551760 0 0 $X=743158 $Y=1551358
X203 2304 1 39 2620 3 2690 OAI21XL $T=944460 1571920 1 0 $X=944458 $Y=1566480
X204 90 1 139 2845 3 2803 OAI21XL $T=990660 1571920 1 0 $X=990658 $Y=1566480
X205 3437 1 3474 3476 3 3424 OAI21XL $T=1148400 1450960 0 0 $X=1148398 $Y=1450558
X206 219 1 161 3498 3 3474 OAI21XL $T=1157640 1450960 0 0 $X=1157638 $Y=1450558
X207 221 1 156 3477 3 3531 OAI21XL $T=1162920 1440880 1 0 $X=1162918 $Y=1435440
X208 3752 1 3764 3729 3 3748 OAI21XL $T=1221660 1461040 0 0 $X=1221658 $Y=1460638
X209 267 1 266 3772 3 3764 OAI21XL $T=1222980 1450960 1 0 $X=1222978 $Y=1445520
X210 4368 1 4417 4353 3 4354 OAI21XL $T=1377420 1571920 0 180 $X=1374780 $Y=1566480
X211 4522 1 4509 4506 3 4491 OAI21XL $T=1411740 1561840 1 180 $X=1409100 $Y=1561438
X212 4506 1 4560 4581 3 4591 OAI21XL $T=1433520 1561840 0 0 $X=1433518 $Y=1561438
X213 4784 1 4725 4726 3 4799 OAI21XL $T=1479720 1481200 1 0 $X=1479718 $Y=1475760
X214 5162 1 399 5071 3 5133 OAI21XL $T=1575420 1551760 1 180 $X=1572780 $Y=1551358
X215 5133 1 5197 5200 3 5204 OAI21XL $T=1574100 1511440 0 0 $X=1574098 $Y=1511038
X216 5200 1 5103 5063 3 5318 OAI21XL $T=1584000 1471120 0 0 $X=1583998 $Y=1470718
X217 404 1 5281 5271 3 5260 OAI21XL $T=1605120 1531600 1 180 $X=1602480 $Y=1531198
X218 5315 1 429 5274 3 430 OAI21XL $T=1618320 1602160 1 0 $X=1618318 $Y=1596720
X219 5465 1 4096 404 3 5421 OAI21XL $T=1636800 1501360 1 180 $X=1634160 $Y=1500958
X220 382 1 5509 4531 3 5460 OAI21XL $T=1658580 1450960 1 180 $X=1655940 $Y=1450558
X221 5521 1 5535 4531 3 5544 OAI21XL $T=1665180 1450960 1 180 $X=1662540 $Y=1450558
X222 313 1 5535 5574 3 5600 OAI21XL $T=1670460 1511440 1 0 $X=1670458 $Y=1506000
X223 439 1 5535 436 3 5574 OAI21XL $T=1673100 1501360 1 0 $X=1673098 $Y=1495920
X224 444 1 5497 453 3 5697 OAI21XL $T=1694220 1440880 0 0 $X=1694218 $Y=1440478
X225 6014 1 467 6016 3 6120 OAI21XL $T=1797180 1511440 1 0 $X=1797178 $Y=1506000
X226 6030 1 6099 6086 3 6117 OAI21XL $T=1807740 1521520 1 0 $X=1807738 $Y=1516080
X227 6121 1 483 6085 3 6099 OAI21XL $T=1813020 1521520 0 0 $X=1813018 $Y=1521118
X228 6097 1 504 6125 3 6206 OAI21XL $T=1814340 1501360 0 0 $X=1814338 $Y=1500958
X229 6204 1 6206 6140 3 6216 OAI21XL $T=1836120 1501360 1 0 $X=1836118 $Y=1495920
X230 6230 1 524 6289 3 6226 OAI21XL $T=1843380 1461040 1 180 $X=1840740 $Y=1460638
X231 6285 1 6306 6304 3 6227 OAI21XL $T=1859220 1481200 0 180 $X=1856580 $Y=1475760
X232 6355 1 6157 6361 3 6285 OAI21XL $T=1870440 1471120 1 0 $X=1870438 $Y=1465680
X233 6414 1 553 6424 3 552 OAI21XL $T=1896840 1450960 0 0 $X=1896838 $Y=1450558
X234 7132 1 614 613 3 7166 OAI21XL $T=2084940 1430800 0 0 $X=2084938 $Y=1430398
X235 7154 1 7138 7132 3 7133 OAI21XL $T=2087580 1450960 1 180 $X=2084940 $Y=1450558
X236 7237 1 7153 7168 3 7169 OAI21XL $T=2096820 1501360 0 180 $X=2094180 $Y=1495920
X237 649 1 653 7736 3 7714 OAI21XL $T=2226180 1602160 1 180 $X=2223540 $Y=1601758
X238 7804 1 7736 7790 3 7795 OAI21XL $T=2242020 1582000 1 180 $X=2239380 $Y=1581598
X239 7766 1 7893 7894 3 7879 OAI21XL $T=2259180 1461040 1 0 $X=2259178 $Y=1455600
X240 669 1 7979 668 3 7957 OAI21XL $T=2287560 1612240 0 180 $X=2284920 $Y=1606800
X241 7997 1 7979 8006 3 7982 OAI21XL $T=2294160 1592080 0 0 $X=2294158 $Y=1591678
X242 8050 1 8006 8068 3 8067 OAI21XL $T=2307360 1582000 0 0 $X=2307358 $Y=1581598
X243 8089 1 8144 8121 3 8154 OAI21XL $T=2331120 1511440 0 0 $X=2331118 $Y=1511038
X244 8086 1 8208 8229 3 8278 OAI21XL $T=2349600 1501360 0 0 $X=2349598 $Y=1500958
X245 8228 1 8166 8199 3 8259 OAI21XL $T=2360820 1491280 1 0 $X=2360818 $Y=1485840
X246 8199 1 8265 8275 3 8230 OAI21XL $T=2366100 1511440 1 0 $X=2366098 $Y=1506000
X247 8351 1 695 8347 3 8326 OAI21XL $T=2384580 1461040 1 180 $X=2381940 $Y=1460638
X248 8423 1 695 8427 3 701 OAI21XL $T=2401740 1430800 0 0 $X=2401738 $Y=1430398
X249 8347 1 8421 8428 3 8440 OAI21XL $T=2404380 1461040 0 0 $X=2404378 $Y=1460638
X250 8510 1 695 8486 3 704 OAI21XL $T=2428800 1440880 1 0 $X=2428798 $Y=1435440
X251 8478 1 8561 8558 3 8562 OAI21XL $T=2444640 1471120 0 0 $X=2444638 $Y=1470718
X252 703 1 575 710 3 8828 OAI21XL $T=2507340 1602160 1 0 $X=2507338 $Y=1596720
X253 726 1 8832 8828 3 728 OAI21XL $T=2516580 1602160 0 180 $X=2513940 $Y=1596720
X254 731 1 8857 8882 3 8804 OAI21XL $T=2523180 1440880 1 0 $X=2523178 $Y=1435440
X255 8780 1 8832 597 3 8979 OAI21XL $T=2541660 1582000 1 0 $X=2541658 $Y=1576560
X256 703 1 594 8979 3 734 OAI21XL $T=2541660 1602160 1 0 $X=2541658 $Y=1596720
X257 717 1 9080 738 3 755 OAI21XL $T=2567400 1612240 1 0 $X=2567398 $Y=1606800
X258 577 1 715 575 3 9188 OAI21XL $T=2597760 1592080 0 0 $X=2597758 $Y=1591678
X259 9187 1 598 9237 3 750 OAI21XL $T=2604360 1561840 0 0 $X=2604358 $Y=1561438
X260 9187 1 9171 717 3 9254 OAI21XL $T=2612280 1561840 1 0 $X=2612278 $Y=1556400
X261 717 1 9270 9254 3 779 OAI21XL $T=2617560 1582000 1 0 $X=2617558 $Y=1576560
X262 28 1566 54 1 3 XOR2X4 $T=662640 1430800 0 0 $X=662638 $Y=1430398
X263 1605 1623 1687 1 3 XOR2X4 $T=678480 1450960 1 0 $X=678478 $Y=1445520
X264 1738 57 55 1 3 XOR2X4 $T=708840 1450960 0 180 $X=697620 $Y=1445520
X265 1844 1804 1929 1 3 XOR2X4 $T=733920 1481200 0 0 $X=733918 $Y=1480798
X266 2472 2496 2604 1 3 XOR2X4 $T=900240 1561840 1 0 $X=900238 $Y=1556400
X267 2546 2446 2577 1 3 XOR2X4 $T=921360 1491280 0 0 $X=921358 $Y=1490878
X268 106 4287 337 1 3 XOR2X4 $T=1345740 1491280 0 0 $X=1345738 $Y=1490878
X269 6660 6615 570 1 3 XOR2X4 $T=1953600 1471120 0 180 $X=1942380 $Y=1465680
X270 6768 6760 583 1 3 XOR2X4 $T=1988580 1450960 0 180 $X=1977360 $Y=1445520
X271 6912 6878 593 1 3 XOR2X4 $T=2012340 1450960 1 180 $X=2001120 $Y=1450558
X272 533 6942 607 1 3 XOR2X4 $T=2019600 1521520 0 0 $X=2019598 $Y=1521118
X273 554 596 608 1 3 XOR2X4 $T=2019600 1551760 1 0 $X=2019598 $Y=1546320
X274 6960 6945 599 1 3 XOR2X4 $T=2036100 1450960 0 180 $X=2024880 $Y=1445520
X275 7709 7685 6779 1 3 XOR2X4 $T=2217600 1561840 1 180 $X=2206380 $Y=1561438
X276 7726 7708 6705 1 3 XOR2X4 $T=2222880 1551760 0 180 $X=2211660 $Y=1546320
X277 8993 8990 8931 1 3 XOR2X4 $T=2564100 1561840 0 180 $X=2552880 $Y=1556400
X278 42 1 3 1651 INVX1 $T=694980 1511440 1 180 $X=693660 $Y=1511038
X279 56 1 3 1636 INVX1 $T=700920 1521520 1 0 $X=700918 $Y=1516080
X280 1722 1 3 1764 INVX1 $T=703560 1481200 0 0 $X=703558 $Y=1480798
X281 1669 1 3 1735 INVX1 $T=703560 1501360 1 0 $X=703558 $Y=1495920
X282 1818 1 3 1803 INVX1 $T=727320 1450960 1 180 $X=726000 $Y=1450558
X283 1840 1 3 1802 INVX1 $T=733260 1602160 1 180 $X=731940 $Y=1601758
X284 80 1 3 88 INVX1 $T=815760 1521520 0 180 $X=814440 $Y=1516080
X285 99 1 3 93 INVX1 $T=825000 1481200 1 180 $X=823680 $Y=1480798
X286 2479 1 3 2480 INVX1 $T=904860 1602160 0 0 $X=904858 $Y=1601758
X287 2477 1 3 2545 INVX1 $T=918060 1450960 1 0 $X=918058 $Y=1445520
X288 2515 1 3 2538 INVX1 $T=920040 1471120 0 0 $X=920038 $Y=1470718
X289 2550 1 3 120 INVX1 $T=933900 1440880 1 0 $X=933898 $Y=1435440
X290 2707 1 3 2704 INVX1 $T=958320 1471120 1 180 $X=957000 $Y=1470718
X291 2724 1 3 2688 INVX1 $T=960960 1521520 0 180 $X=959640 $Y=1516080
X292 2790 1 3 2686 INVX1 $T=979440 1511440 1 180 $X=978120 $Y=1511038
X293 2803 1 3 2809 INVX1 $T=980760 1551760 0 0 $X=980758 $Y=1551358
X294 2826 1 3 2789 INVX1 $T=984720 1481200 1 180 $X=983400 $Y=1480798
X295 31 1 3 2689 INVX1 $T=993960 1571920 0 0 $X=993958 $Y=1571518
X296 2907 1 3 2903 INVX1 $T=1001880 1481200 0 180 $X=1000560 $Y=1475760
X297 2918 1 3 2949 INVX1 $T=1007160 1491280 0 0 $X=1007158 $Y=1490878
X298 153 1 3 147 INVX1 $T=1027620 1461040 0 0 $X=1027618 $Y=1460638
X299 3111 1 3 2948 INVX1 $T=1044780 1521520 1 180 $X=1043460 $Y=1521118
X300 36 1 3 2905 INVX1 $T=1047420 1582000 0 180 $X=1046100 $Y=1576560
X301 2973 1 3 3052 INVX1 $T=1055340 1501360 0 180 $X=1054020 $Y=1495920
X302 177 1 3 3159 INVX1 $T=1072500 1491280 0 0 $X=1072498 $Y=1490878
X303 3158 1 3 3171 INVX1 $T=1075140 1481200 1 0 $X=1075138 $Y=1475760
X304 3177 1 3 180 INVX1 $T=1079100 1450960 0 180 $X=1077780 $Y=1445520
X305 130 1 3 3261 INVX1 $T=1098240 1592080 1 0 $X=1098238 $Y=1586640
X306 3292 1 3 3231 INVX1 $T=1102200 1481200 1 180 $X=1100880 $Y=1480798
X307 39 1 3 196 INVX1 $T=1135200 1612240 0 0 $X=1135198 $Y=1611838
X308 195 1 3 3435 INVX1 $T=1143120 1440880 1 0 $X=1143118 $Y=1435440
X309 201 1 3 3481 INVX1 $T=1153680 1471120 1 0 $X=1153678 $Y=1465680
X310 99 1 3 3493 INVX1 $T=1155660 1571920 1 0 $X=1155658 $Y=1566480
X311 203 1 3 236 INVX1 $T=1182060 1511440 0 0 $X=1182058 $Y=1511038
X312 253 1 3 257 INVX1 $T=1205160 1430800 0 0 $X=1205158 $Y=1430398
X313 285 1 3 262 INVX1 $T=1215060 1430800 1 180 $X=1213740 $Y=1430398
X314 274 1 3 3796 INVX1 $T=1228920 1471120 0 0 $X=1228918 $Y=1470718
X315 296 1 3 286 INVX1 $T=1259280 1440880 0 180 $X=1257960 $Y=1435440
X316 4040 1 3 4056 INVX1 $T=1298220 1491280 0 0 $X=1298218 $Y=1490878
X317 4057 1 3 4061 INVX1 $T=1298880 1571920 0 0 $X=1298878 $Y=1571518
X318 4097 1 3 4112 INVX1 $T=1310100 1551760 1 0 $X=1310098 $Y=1546320
X319 4101 1 3 4145 INVX1 $T=1315380 1501360 0 0 $X=1315378 $Y=1500958
X320 328 1 3 4146 INVX1 $T=1330560 1571920 0 180 $X=1329240 $Y=1566480
X321 341 1 3 160 INVX1 $T=1364220 1461040 0 180 $X=1362900 $Y=1455600
X322 343 1 3 4417 INVX1 $T=1393920 1571920 1 0 $X=1393918 $Y=1566480
X323 345 1 3 4416 INVX1 $T=1395900 1501360 0 180 $X=1394580 $Y=1495920
X324 4394 1 3 4476 INVX1 $T=1399200 1491280 0 0 $X=1399198 $Y=1490878
X325 350 1 3 4479 INVX1 $T=1405800 1531600 0 180 $X=1404480 $Y=1526160
X326 4507 1 3 4477 INVX1 $T=1413720 1511440 0 180 $X=1412400 $Y=1506000
X327 4486 1 3 4527 INVX1 $T=1417020 1501360 1 0 $X=1417018 $Y=1495920
X328 4550 1 3 4509 INVX1 $T=1427580 1571920 1 0 $X=1427578 $Y=1566480
X329 4585 1 3 4598 INVX1 $T=1435500 1511440 1 0 $X=1435498 $Y=1506000
X330 359 1 3 4727 INVX1 $T=1469160 1531600 1 0 $X=1469158 $Y=1526160
X331 371 1 3 4851 INVX1 $T=1497540 1551760 1 0 $X=1497538 $Y=1546320
X332 4041 1 3 387 INVX1 $T=1519320 1531600 0 0 $X=1519318 $Y=1531198
X333 4227 1 3 4096 INVX1 $T=1523280 1521520 1 180 $X=1521960 $Y=1521118
X334 391 1 3 5038 INVX1 $T=1537800 1551760 0 0 $X=1537798 $Y=1551358
X335 5046 1 3 5070 INVX1 $T=1545720 1501360 0 0 $X=1545718 $Y=1500958
X336 5025 1 3 5022 INVX1 $T=1551000 1521520 1 0 $X=1550998 $Y=1516080
X337 5225 1 3 5110 INVX1 $T=1565520 1501360 1 180 $X=1564200 $Y=1500958
X338 5063 1 3 5180 INVX1 $T=1572120 1531600 1 0 $X=1572118 $Y=1526160
X339 4748 1 3 5199 INVX1 $T=1574100 1450960 0 0 $X=1574098 $Y=1450558
X340 5158 1 3 4744 INVX1 $T=1575420 1582000 1 180 $X=1574100 $Y=1581598
X341 5237 1 3 5201 INVX1 $T=1584660 1582000 1 0 $X=1584658 $Y=1576560
X342 417 1 3 418 INVX1 $T=1589940 1430800 0 0 $X=1589938 $Y=1430398
X343 5271 1 3 5153 INVX1 $T=1595220 1531600 1 0 $X=1595218 $Y=1526160
X344 5281 1 3 5194 INVX1 $T=1597860 1541680 1 0 $X=1597858 $Y=1536240
X345 399 1 3 420 INVX1 $T=1597860 1602160 1 0 $X=1597858 $Y=1596720
X346 5321 1 3 5197 INVX1 $T=1607100 1521520 1 180 $X=1605780 $Y=1521118
X347 404 1 3 416 INVX1 $T=1608420 1541680 1 0 $X=1608418 $Y=1536240
X348 5326 1 3 5324 INVX1 $T=1608420 1582000 0 0 $X=1608418 $Y=1581598
X349 5327 1 3 5259 INVX1 $T=1609740 1511440 1 180 $X=1608420 $Y=1511038
X350 5103 1 3 5253 INVX1 $T=1611060 1491280 1 0 $X=1611058 $Y=1485840
X351 424 1 3 5355 INVX1 $T=1616340 1582000 1 0 $X=1616338 $Y=1576560
X352 5274 1 3 5129 INVX1 $T=1617660 1561840 0 180 $X=1616340 $Y=1556400
X353 5380 1 3 5352 INVX1 $T=1623600 1571920 1 0 $X=1623598 $Y=1566480
X354 5269 1 3 5388 INVX1 $T=1625580 1501360 0 180 $X=1624260 $Y=1495920
X355 5361 1 3 5298 INVX1 $T=1625580 1551760 1 180 $X=1624260 $Y=1551358
X356 5431 1 3 5391 INVX1 $T=1634820 1491280 0 180 $X=1633500 $Y=1485840
X357 5352 1 3 5419 INVX1 $T=1634160 1531600 1 0 $X=1634158 $Y=1526160
X358 5390 1 3 5399 INVX1 $T=1634820 1592080 1 0 $X=1634818 $Y=1586640
X359 5254 1 3 5150 INVX1 $T=1640760 1521520 0 0 $X=1640758 $Y=1521118
X360 5220 1 3 5198 INVX1 $T=1644060 1571920 1 180 $X=1642740 $Y=1571518
X361 5246 1 3 5497 INVX1 $T=1650000 1440880 0 0 $X=1649998 $Y=1440478
X362 4531 1 3 439 INVX1 $T=1655280 1450960 1 0 $X=1655278 $Y=1445520
X363 5509 1 3 5498 INVX1 $T=1656600 1511440 0 180 $X=1655280 $Y=1506000
X364 440 1 3 5494 INVX1 $T=1659240 1471120 1 180 $X=1657920 $Y=1470718
X365 5533 1 3 5535 INVX1 $T=1661220 1450960 0 180 $X=1659900 $Y=1445520
X366 5535 1 3 5524 INVX1 $T=1661880 1511440 0 180 $X=1660560 $Y=1506000
X367 5523 1 3 5236 INVX1 $T=1663200 1471120 1 180 $X=1661880 $Y=1470718
X368 377 1 3 5560 INVX1 $T=1667820 1612240 0 0 $X=1667818 $Y=1611838
X369 450 1 3 5577 INVX1 $T=1690920 1481200 0 180 $X=1689600 $Y=1475760
X370 415 1 3 427 INVX1 $T=1705440 1571920 0 0 $X=1705438 $Y=1571518
X371 419 1 3 5465 INVX1 $T=1708080 1501360 0 0 $X=1708078 $Y=1500958
X372 469 1 3 5897 INVX1 $T=1752960 1491280 1 0 $X=1752958 $Y=1485840
X373 5698 1 3 5952 INVX1 $T=1763520 1491280 0 0 $X=1763518 $Y=1490878
X374 398 1 3 414 INVX1 $T=1765500 1592080 1 0 $X=1765498 $Y=1586640
X375 475 1 3 5968 INVX1 $T=1772100 1501360 1 0 $X=1772098 $Y=1495920
X376 479 1 3 6014 INVX1 $T=1781340 1511440 1 0 $X=1781338 $Y=1506000
X377 468 1 3 482 INVX1 $T=1785300 1430800 0 0 $X=1785298 $Y=1430398
X378 481 1 3 6048 INVX1 $T=1785960 1521520 0 0 $X=1785958 $Y=1521118
X379 486 1 3 6018 INVX1 $T=1788600 1521520 1 0 $X=1788598 $Y=1516080
X380 496 1 3 6097 INVX1 $T=1804440 1501360 1 0 $X=1804438 $Y=1495920
X381 473 1 3 6100 INVX1 $T=1807080 1491280 1 0 $X=1807078 $Y=1485840
X382 499 1 3 6121 INVX1 $T=1809720 1531600 0 0 $X=1809718 $Y=1531198
X383 513 1 3 6207 INVX1 $T=1825560 1521520 0 0 $X=1825558 $Y=1521118
X384 524 1 3 477 INVX1 $T=1827540 1612240 1 180 $X=1826220 $Y=1611838
X385 6187 1 3 6178 INVX1 $T=1834800 1551760 1 180 $X=1833480 $Y=1551358
X386 523 1 3 6231 INVX1 $T=1838760 1521520 0 0 $X=1838758 $Y=1521118
X387 468 1 3 6230 INVX1 $T=1841400 1450960 1 0 $X=1841398 $Y=1445520
X388 6227 1 3 6233 INVX1 $T=1841400 1481200 1 0 $X=1841398 $Y=1475760
X389 506 1 3 478 INVX1 $T=1848660 1561840 1 0 $X=1848658 $Y=1556400
X390 489 1 3 6302 INVX1 $T=1854600 1450960 1 0 $X=1854598 $Y=1445520
X391 558 1 3 518 INVX1 $T=1855920 1582000 1 180 $X=1854600 $Y=1581598
X392 6326 1 3 6324 INVX1 $T=1863180 1511440 1 180 $X=1861860 $Y=1511038
X393 534 1 3 514 INVX1 $T=1863180 1551760 1 180 $X=1861860 $Y=1551358
X394 535 1 3 6364 INVX1 $T=1867140 1501360 0 0 $X=1867138 $Y=1500958
X395 509 1 3 6355 INVX1 $T=1869780 1450960 0 0 $X=1869778 $Y=1450558
X396 509 1 3 6414 INVX1 $T=1872420 1440880 0 0 $X=1872418 $Y=1440478
X397 549 1 3 6157 INVX1 $T=1886940 1592080 1 180 $X=1885620 $Y=1591678
X398 551 1 3 6422 INVX1 $T=1890900 1440880 0 0 $X=1890898 $Y=1440478
X399 551 1 3 6346 INVX1 $T=1893540 1471120 1 0 $X=1893538 $Y=1465680
X400 556 1 3 6398 INVX1 $T=1901460 1440880 1 0 $X=1901458 $Y=1435440
X401 6495 1 3 506 INVX1 $T=1907400 1551760 0 180 $X=1906080 $Y=1546320
X402 553 1 3 520 INVX1 $T=1944360 1450960 0 180 $X=1943040 $Y=1445520
X403 6686 1 3 6664 INVX1 $T=1960200 1450960 0 0 $X=1960198 $Y=1450558
X404 586 1 3 6795 INVX1 $T=1987260 1551760 1 0 $X=1987258 $Y=1546320
X405 591 1 3 6800 INVX1 $T=1997160 1561840 1 180 $X=1995840 $Y=1561438
X406 6878 1 3 6900 INVX1 $T=2013660 1491280 0 0 $X=2013658 $Y=1490878
X407 7050 1 3 7068 INVX1 $T=2064480 1501360 1 0 $X=2064478 $Y=1495920
X408 7100 1 3 7109 INVX1 $T=2073720 1511440 0 0 $X=2073718 $Y=1511038
X409 7169 1 3 7138 INVX1 $T=2094840 1461040 1 0 $X=2094838 $Y=1455600
X410 7171 1 3 7221 INVX1 $T=2094840 1582000 1 0 $X=2094838 $Y=1576560
X411 7253 1 3 7369 INVX1 $T=2141700 1571920 1 0 $X=2141698 $Y=1566480
X412 637 1 3 632 INVX1 $T=2153580 1612240 1 180 $X=2152260 $Y=1611838
X413 7488 1 3 7425 INVX1 $T=2170740 1571920 1 180 $X=2169420 $Y=1571518
X414 7511 1 3 7359 INVX1 $T=2172060 1481200 1 180 $X=2170740 $Y=1480798
X415 7512 1 3 7474 INVX1 $T=2174700 1561840 0 180 $X=2173380 $Y=1556400
X416 7473 1 3 643 INVX1 $T=2176020 1430800 0 0 $X=2176018 $Y=1430398
X417 644 1 3 7548 INVX1 $T=2185260 1582000 1 180 $X=2183940 $Y=1581598
X418 7442 1 3 7526 INVX1 $T=2187900 1521520 1 180 $X=2186580 $Y=1521118
X419 7571 1 3 7587 INVX1 $T=2190540 1461040 1 0 $X=2190538 $Y=1455600
X420 7652 1 3 7557 INVX1 $T=2202420 1541680 0 180 $X=2201100 $Y=1536240
X421 7608 1 3 7651 INVX1 $T=2209680 1491280 1 180 $X=2208360 $Y=1490878
X422 651 1 3 7686 INVX1 $T=2213640 1592080 1 180 $X=2212320 $Y=1591678
X423 7757 1 3 7735 INVX1 $T=2232120 1582000 0 180 $X=2230800 $Y=1576560
X424 7772 1 3 7732 INVX1 $T=2234100 1582000 1 0 $X=2234098 $Y=1576560
X425 7683 1 3 7754 INVX1 $T=2238720 1461040 0 0 $X=2238718 $Y=1460638
X426 657 1 3 7647 INVX1 $T=2240040 1602160 1 180 $X=2238720 $Y=1601758
X427 7880 1 3 7789 INVX1 $T=2258520 1582000 0 180 $X=2257200 $Y=1576560
X428 7825 1 3 7865 INVX1 $T=2259180 1541680 0 180 $X=2257860 $Y=1536240
X429 7810 1 3 7878 INVX1 $T=2262480 1541680 1 180 $X=2261160 $Y=1541278
X430 7882 1 3 7897 INVX1 $T=2269080 1531600 0 180 $X=2267760 $Y=1526160
X431 7933 1 3 7649 INVX1 $T=2274360 1481200 0 180 $X=2273040 $Y=1475760
X432 7972 1 3 7914 INVX1 $T=2281620 1541680 0 180 $X=2280300 $Y=1536240
X433 7960 1 3 7788 INVX1 $T=2282280 1471120 1 180 $X=2280960 $Y=1470718
X434 667 1 3 7979 INVX1 $T=2282940 1592080 0 0 $X=2282938 $Y=1591678
X435 8063 1 3 7670 INVX1 $T=2293500 1481200 0 180 $X=2292180 $Y=1475760
X436 668 1 3 8065 INVX1 $T=2301420 1602160 0 0 $X=2301418 $Y=1601758
X437 8088 1 3 7913 INVX1 $T=2313300 1471120 1 180 $X=2311980 $Y=1470718
X438 8086 1 3 8064 INVX1 $T=2319240 1501360 0 0 $X=2319238 $Y=1500958
X439 675 1 3 8069 INVX1 $T=2322540 1612240 0 0 $X=2322538 $Y=1611838
X440 8134 1 3 8117 INVX1 $T=2329140 1440880 0 180 $X=2327820 $Y=1435440
X441 685 1 3 8115 INVX1 $T=2344980 1440880 1 180 $X=2343660 $Y=1440478
X442 8235 1 3 8207 INVX1 $T=2354880 1461040 0 180 $X=2353560 $Y=1455600
X443 598 1 3 6661 INVX1 $T=2355540 1612240 1 0 $X=2355538 $Y=1606800
X444 8334 1 3 8244 INVX1 $T=2384580 1450960 1 0 $X=2384578 $Y=1445520
X445 8424 1 3 8423 INVX1 $T=2402400 1440880 0 180 $X=2401080 $Y=1435440
X446 677 1 3 8374 INVX1 $T=2402400 1592080 1 180 $X=2401080 $Y=1591678
X447 575 1 3 6695 INVX1 $T=2421540 1582000 1 0 $X=2421538 $Y=1576560
X448 8901 1 3 7810 INVX1 $T=2495460 1551760 1 180 $X=2494140 $Y=1551358
X449 598 1 3 717 INVX1 $T=2507340 1571920 1 0 $X=2507338 $Y=1566480
X450 594 1 3 8780 INVX1 $T=2515920 1582000 1 0 $X=2515918 $Y=1576560
X451 575 1 3 726 INVX1 $T=2526480 1571920 0 0 $X=2526478 $Y=1571518
X452 703 1 3 8832 INVX1 $T=2531100 1602160 1 0 $X=2531098 $Y=1596720
X453 752 1 3 754 INVX1 $T=2607660 1430800 0 0 $X=2607658 $Y=1430398
X454 9171 1 3 9237 INVX1 $T=2608980 1561840 0 180 $X=2607660 $Y=1556400
X455 1565 1562 3 29 1566 1 AOI21X2 $T=668580 1461040 1 180 $X=663960 $Y=1460638
X456 1565 1560 3 51 1623 1 AOI21X2 $T=687060 1461040 0 180 $X=682440 $Y=1455600
X457 1565 1764 3 1801 1804 1 AOI21X2 $T=721380 1481200 0 0 $X=721378 $Y=1480798
X458 1850 1823 3 1826 1839 1 AOI21X2 $T=733920 1571920 1 180 $X=729300 $Y=1571518
X459 112 115 3 2480 2478 1 AOI21X2 $T=908820 1602160 0 180 $X=904200 $Y=1596720
X460 2533 2538 3 2545 2509 1 AOI21X2 $T=920040 1450960 0 0 $X=920038 $Y=1450558
X461 2446 2534 3 2538 119 1 AOI21X2 $T=925980 1471120 0 180 $X=921360 $Y=1465680
X462 2772 2762 3 2789 2727 1 AOI21X2 $T=974820 1481200 0 0 $X=974818 $Y=1480798
X463 3018 163 3 3008 162 1 AOI21X2 $T=1036200 1501360 0 180 $X=1031580 $Y=1495920
X464 4477 4414 3 4476 4489 1 AOI21X2 $T=1409100 1491280 1 180 $X=1404480 $Y=1490878
X465 4582 4550 3 4591 4599 1 AOI21X2 $T=1434840 1571920 1 0 $X=1434838 $Y=1566480
X466 6757 584 3 6795 6799 1 AOI21X2 $T=1985940 1541680 1 0 $X=1985938 $Y=1536240
X467 6762 6795 3 6800 6761 1 AOI21X2 $T=1989240 1551760 0 0 $X=1989238 $Y=1551358
X468 7167 7169 3 7166 617 1 AOI21X2 $T=2094180 1430800 0 0 $X=2094178 $Y=1430398
X469 618 7222 3 7221 7253 1 AOI21X2 $T=2102760 1582000 1 0 $X=2102758 $Y=1576560
X470 7687 651 3 7714 7708 1 AOI21X2 $T=2214960 1602160 0 0 $X=2214958 $Y=1601758
X471 7856 7861 3 7897 7896 1 AOI21X2 $T=2259180 1531600 1 0 $X=2259178 $Y=1526160
X472 7897 7862 3 7914 7825 1 AOI21X2 $T=2264460 1541680 1 0 $X=2264458 $Y=1536240
X473 676 8115 3 8117 8066 1 AOI21X2 $T=2319240 1440880 1 0 $X=2319238 $Y=1435440
X474 9095 9086 3 9082 8990 1 AOI21X2 $T=2572680 1551760 1 180 $X=2568060 $Y=1551358
X475 3 1598 1581 43 1 NOR2X1 $T=675840 1531600 0 0 $X=675838 $Y=1531198
X476 3 1872 1818 69 1 NOR2X1 $T=733920 1450960 1 180 $X=731940 $Y=1450558
X477 3 64 1840 1817 1 NOR2X1 $T=732600 1612240 0 0 $X=732598 $Y=1611838
X478 3 1878 1856 1818 1 NOR2X1 $T=739200 1461040 0 180 $X=737220 $Y=1455600
X479 3 1997 1927 1872 1 NOR2X1 $T=752400 1450960 1 180 $X=750420 $Y=1450558
X480 3 1928 1930 1819 1 NOR2X1 $T=756360 1561840 0 0 $X=756358 $Y=1561438
X481 3 2781 2790 2765 1 NOR2X1 $T=976800 1501360 0 0 $X=976798 $Y=1500958
X482 3 2837 2819 2833 1 NOR2X1 $T=989340 1602160 0 180 $X=987360 $Y=1596720
X483 3 144 146 2790 1 NOR2X1 $T=1003200 1511440 1 180 $X=1001220 $Y=1511038
X484 3 155 148 2837 1 NOR2X1 $T=1013760 1612240 0 180 $X=1011780 $Y=1606800
X485 3 3038 2907 3031 1 NOR2X1 $T=1032900 1481200 0 0 $X=1032898 $Y=1480798
X486 3 153 174 3111 1 NOR2X1 $T=1060620 1551760 0 180 $X=1058640 $Y=1546320
X487 3 4368 4305 4350 1 NOR2X1 $T=1372800 1561840 1 180 $X=1370820 $Y=1561438
X488 3 4490 4488 4522 1 NOR2X1 $T=1415040 1571920 1 0 $X=1415038 $Y=1566480
X489 3 354 353 4524 1 NOR2X1 $T=1421640 1612240 0 180 $X=1419660 $Y=1606800
X490 3 4522 4560 4582 1 NOR2X1 $T=1426260 1561840 0 0 $X=1426258 $Y=1561438
X491 3 4293 4590 4577 1 NOR2X1 $T=1435500 1471120 0 0 $X=1435498 $Y=1470718
X492 3 4597 357 4635 1 NOR2X1 $T=1446060 1430800 0 0 $X=1446058 $Y=1430398
X493 3 4532 4637 4585 1 NOR2X1 $T=1446720 1511440 0 0 $X=1446718 $Y=1511038
X494 3 358 355 4683 1 NOR2X1 $T=1451340 1481200 0 180 $X=1449360 $Y=1475760
X495 3 4292 4693 4692 1 NOR2X1 $T=1453980 1461040 1 0 $X=1453978 $Y=1455600
X496 3 364 361 4779 1 NOR2X1 $T=1472460 1541680 0 0 $X=1472458 $Y=1541278
X497 3 4770 365 4704 1 NOR2X1 $T=1475100 1430800 1 180 $X=1473120 $Y=1430398
X498 3 4583 4785 4784 1 NOR2X1 $T=1479720 1491280 1 0 $X=1479718 $Y=1485840
X499 3 4205 4817 4870 1 NOR2X1 $T=1490280 1450960 1 0 $X=1490278 $Y=1445520
X500 3 5025 5063 5050 1 NOR2X1 $T=1549680 1531600 0 180 $X=1547700 $Y=1526160
X501 3 5153 5150 5158 1 NOR2X1 $T=1563540 1541680 0 0 $X=1563538 $Y=1541278
X502 3 5063 5195 328 1 NOR2X1 $T=1573440 1521520 1 0 $X=1573438 $Y=1516080
X503 3 5158 387 5237 1 NOR2X1 $T=1582020 1592080 1 0 $X=1582018 $Y=1586640
X504 3 5063 5200 5254 1 NOR2X1 $T=1584660 1521520 1 0 $X=1584658 $Y=1516080
X505 3 5025 5253 5271 1 NOR2X1 $T=1589940 1521520 1 0 $X=1589938 $Y=1516080
X506 3 5200 5180 5281 1 NOR2X1 $T=1595220 1521520 0 0 $X=1595218 $Y=1521118
X507 3 420 5256 5218 1 NOR2X1 $T=1595220 1582000 0 0 $X=1595218 $Y=1581598
X508 3 328 403 5247 1 NOR2X1 $T=1597200 1582000 0 180 $X=1595220 $Y=1576560
X509 3 419 4745 5516 1 NOR2X1 $T=1681020 1582000 1 0 $X=1681018 $Y=1576560
X510 3 442 5539 454 1 NOR2X1 $T=1691580 1450960 1 0 $X=1691578 $Y=1445520
X511 3 5352 4723 5775 1 NOR2X1 $T=1725900 1571920 0 0 $X=1725898 $Y=1571518
X512 3 5968 5952 5950 1 NOR2X1 $T=1772760 1491280 1 180 $X=1770780 $Y=1490878
X513 3 502 6039 6156 1 NOR2X1 $T=1812360 1450960 1 0 $X=1812358 $Y=1445520
X514 3 6191 6190 6159 1 NOR2X1 $T=1832160 1450960 0 180 $X=1830180 $Y=1445520
X515 3 518 510 6292 1 NOR2X1 $T=1853940 1592080 1 0 $X=1853938 $Y=1586640
X516 3 531 483 565 1 NOR2X1 $T=1931160 1430800 0 0 $X=1931158 $Y=1430398
X517 3 6661 572 6345 1 NOR2X1 $T=1950300 1602160 0 180 $X=1948320 $Y=1596720
X518 3 588 576 6542 1 NOR2X1 $T=1960860 1592080 1 180 $X=1958880 $Y=1591678
X519 3 6930 6946 7012 1 NOR2X1 $T=2046660 1481200 1 0 $X=2046658 $Y=1475760
X520 3 7154 614 7167 1 NOR2X1 $T=2090880 1440880 1 0 $X=2090878 $Y=1435440
X521 3 568 7139 7154 1 NOR2X1 $T=2097480 1450960 1 180 $X=2095500 $Y=1450558
X522 3 571 608 7237 1 NOR2X1 $T=2114640 1501360 0 180 $X=2112660 $Y=1495920
X523 3 629 7342 7331 1 NOR2X1 $T=2137740 1521520 1 180 $X=2135760 $Y=1521118
X524 3 649 7647 7687 1 NOR2X1 $T=2211000 1602160 1 180 $X=2209020 $Y=1601758
X525 3 7788 655 7783 1 NOR2X1 $T=2239380 1461040 0 180 $X=2237400 $Y=1455600
X526 3 7804 649 7813 1 NOR2X1 $T=2242680 1602160 0 180 $X=2240700 $Y=1596720
X527 3 7783 7893 7874 1 NOR2X1 $T=2262480 1450960 0 0 $X=2262478 $Y=1450558
X528 3 673 7990 8050 1 NOR2X1 $T=2298120 1582000 1 180 $X=2296140 $Y=1581598
X529 3 8050 7997 8051 1 NOR2X1 $T=2301420 1592080 1 0 $X=2301418 $Y=1586640
X530 3 8119 8101 8085 1 NOR2X1 $T=2321220 1521520 1 180 $X=2319240 $Y=1521118
X531 3 8085 8144 8137 1 NOR2X1 $T=2332440 1521520 1 0 $X=2332438 $Y=1516080
X532 3 8122 8157 8144 1 NOR2X1 $T=2335740 1541680 1 180 $X=2333760 $Y=1541278
X533 3 8207 687 685 1 NOR2X1 $T=2349600 1450960 1 180 $X=2347620 $Y=1450558
X534 3 8228 8265 8200 1 NOR2X1 $T=2366100 1521520 0 180 $X=2364120 $Y=1516080
X535 3 8247 8245 8228 1 NOR2X1 $T=2367420 1531600 0 180 $X=2365440 $Y=1526160
X536 3 8304 8303 8265 1 NOR2X1 $T=2376660 1521520 1 180 $X=2374680 $Y=1521118
X537 3 8345 8353 8351 1 NOR2X1 $T=2391840 1481200 1 180 $X=2389860 $Y=1480798
X538 3 8421 8351 8424 1 NOR2X1 $T=2400420 1461040 1 0 $X=2400418 $Y=1455600
X539 3 8438 8422 8421 1 NOR2X1 $T=2402400 1501360 0 180 $X=2400420 $Y=1495920
X540 3 8511 8508 8497 1 NOR2X1 $T=2428800 1481200 0 180 $X=2426820 $Y=1475760
X541 3 8561 8497 8560 1 NOR2X1 $T=2443320 1450960 1 180 $X=2441340 $Y=1450558
X542 3 8627 8551 8561 1 NOR2X1 $T=2457180 1481200 0 180 $X=2455200 $Y=1475760
X543 3 8671 8682 713 1 NOR2X1 $T=2478960 1450960 0 0 $X=2478958 $Y=1450558
X544 3 8738 8711 719 1 NOR2X1 $T=2485560 1440880 0 0 $X=2485558 $Y=1440478
X545 3 8857 729 8786 1 NOR2X1 $T=2517900 1430800 1 180 $X=2515920 $Y=1430398
X546 3 8883 8781 729 1 NOR2X1 $T=2519220 1450960 0 180 $X=2517240 $Y=1445520
X547 3 8884 8910 8857 1 NOR2X1 $T=2533080 1450960 0 180 $X=2531100 $Y=1445520
X548 1722 1669 1 3 1560 NOR2X2 $T=693660 1481200 1 180 $X=690360 $Y=1480798
X549 1661 53 1 3 1669 NOR2X2 $T=693000 1531600 1 0 $X=692998 $Y=1526160
X550 1723 59 1 3 1722 NOR2X2 $T=703560 1592080 1 0 $X=703558 $Y=1586640
X551 1819 1849 1 3 1850 NOR2X2 $T=739860 1561840 0 180 $X=736560 $Y=1556400
X552 1959 1960 1 3 1840 NOR2X2 $T=757020 1602160 0 180 $X=753720 $Y=1596720
X553 1992 1993 1 3 1849 NOR2X2 $T=766260 1551760 1 180 $X=762960 $Y=1551358
X554 1961 2347 1 3 2394 NOR2X2 $T=880440 1501360 1 0 $X=880438 $Y=1495920
X555 2394 2395 1 3 2420 NOR2X2 $T=895620 1501360 0 180 $X=892320 $Y=1495920
X556 141 140 1 3 2781 NOR2X2 $T=990660 1521520 0 180 $X=987360 $Y=1516080
X557 152 154 1 3 2819 NOR2X2 $T=1007820 1602160 0 180 $X=1004520 $Y=1596720
X558 2740 342 1 3 4368 NOR2X2 $T=1372140 1612240 1 0 $X=1372138 $Y=1606800
X559 4617 4487 1 3 4560 NOR2X2 $T=1441440 1561840 0 0 $X=1441438 $Y=1561438
X560 3883 358 1 3 3980 NOR2X2 $T=1452660 1531600 1 180 $X=1449360 $Y=1531198
X561 4800 4784 1 3 4812 NOR2X2 $T=1481700 1481200 0 0 $X=1481698 $Y=1480798
X562 4723 5039 1 3 4856 NOR2X2 $T=1517340 1571920 0 180 $X=1514040 $Y=1566480
X563 5131 5101 1 3 5148 NOR2X2 $T=1560900 1501360 0 0 $X=1560898 $Y=1500958
X564 5516 5560 1 3 460 NOR2X2 $T=1681020 1612240 0 0 $X=1681018 $Y=1611838
X565 5894 358 1 3 5896 NOR2X2 $T=1752300 1551760 1 0 $X=1752298 $Y=1546320
X566 5950 5912 1 3 5967 NOR2X2 $T=1769460 1481200 0 0 $X=1769458 $Y=1480798
X567 539 533 1 3 6498 NOR2X2 $T=1912020 1511440 1 180 $X=1908720 $Y=1511038
X568 7307 7312 1 3 7306 NOR2X2 $T=2128500 1521520 0 180 $X=2125200 $Y=1516080
X569 7712 650 1 3 7668 NOR2X2 $T=2213640 1511440 1 180 $X=2210340 $Y=1511038
X570 7794 7711 1 3 7786 NOR2X2 $T=2238720 1491280 0 0 $X=2238718 $Y=1490878
X571 7824 659 1 3 7711 NOR2X2 $T=2244660 1501360 0 180 $X=2241360 $Y=1495920
X572 662 7913 1 3 7893 NOR2X2 $T=2270400 1461040 1 0 $X=2270398 $Y=1455600
X573 670 7991 1 3 666 NOR2X2 $T=2280960 1430800 1 180 $X=2277660 $Y=1430398
X574 694 8244 1 3 684 NOR2X2 $T=2356200 1440880 1 0 $X=2356198 $Y=1435440
X575 1822 72 1 3 1848 OR2XL $T=740520 1521520 0 180 $X=737880 $Y=1516080
X576 108 102 1 3 2196 OR2XL $T=845460 1440880 1 180 $X=842820 $Y=1440478
X577 1961 2347 1 3 2348 OR2XL $T=869880 1501360 1 0 $X=869878 $Y=1495920
X578 159 3481 1 3 3498 OR2XL $T=1165560 1461040 1 180 $X=1162920 $Y=1460638
X579 265 262 1 3 3772 OR2XL $T=1228260 1440880 0 180 $X=1225620 $Y=1435440
X580 4041 174 1 3 4212 OR2XL $T=1337160 1541680 0 0 $X=1337158 $Y=1541278
X581 4227 322 1 3 4249 OR2XL $T=1343760 1541680 1 0 $X=1343758 $Y=1536240
X582 4227 323 1 3 4233 OR2XL $T=1349040 1531600 0 180 $X=1346400 $Y=1526160
X583 4227 245 1 3 4304 OR2XL $T=1359600 1531600 0 180 $X=1356960 $Y=1526160
X584 4041 341 1 3 4302 OR2XL $T=1368840 1521520 1 180 $X=1366200 $Y=1521118
X585 494 6048 1 3 6085 OR2XL $T=1797180 1521520 0 0 $X=1797178 $Y=1521118
X586 498 6100 1 3 6125 OR2XL $T=1809060 1501360 1 0 $X=1809058 $Y=1495920
X587 501 6302 1 3 6289 OR2XL $T=1869120 1461040 1 180 $X=1866480 $Y=1460638
X588 536 6346 1 3 6361 OR2XL $T=1883640 1481200 0 180 $X=1881000 $Y=1475760
X589 550 6422 1 3 6424 OR2XL $T=1890240 1450960 1 0 $X=1890238 $Y=1445520
X590 571 6600 1 3 595 OR2XL $T=2007720 1511440 1 0 $X=2007718 $Y=1506000
X591 571 567 1 3 7119 OR2XL $T=2089560 1521520 0 180 $X=2086920 $Y=1516080
X592 715 710 1 3 8699 OR2XL $T=2485560 1551760 1 180 $X=2482920 $Y=1551358
X593 755 566 1 3 757 OR2XL $T=2612280 1612240 0 0 $X=2612278 $Y=1611838
X594 1560 5 33 1 3 NAND2X2 $T=664620 1440880 0 0 $X=664618 $Y=1440478
X595 114 2478 2427 1 3 NAND2X2 $T=898920 1571920 1 180 $X=895620 $Y=1571518
X596 2772 2765 2770 1 3 NAND2X2 $T=974160 1491280 0 0 $X=974158 $Y=1490878
X597 131 134 2725 1 3 NAND2X2 $T=978120 1440880 0 0 $X=978118 $Y=1440478
X598 146 144 2724 1 3 NAND2X2 $T=999240 1521520 1 0 $X=999238 $Y=1516080
X599 148 155 2834 1 3 NAND2X2 $T=1000560 1612240 1 0 $X=1000558 $Y=1606800
X600 2938 2948 2970 1 3 NAND2X2 $T=1028280 1491280 1 0 $X=1028278 $Y=1485840
X601 2604 336 4289 1 3 NAND2X2 $T=1354320 1561840 0 180 $X=1351020 $Y=1556400
X602 2740 342 4353 1 3 NAND2X2 $T=1368180 1602160 1 180 $X=1364880 $Y=1601758
X603 4414 4478 4486 1 3 NAND2X2 $T=1409100 1501360 0 180 $X=1405800 $Y=1495920
X604 4475 4527 4558 1 3 NAND2X2 $T=1424280 1501360 1 0 $X=1424278 $Y=1495920
X605 4855 4510 4815 1 3 NAND2X2 $T=1496220 1481200 1 0 $X=1496218 $Y=1475760
X606 392 5127 5102 1 3 NAND2X2 $T=1553640 1582000 0 180 $X=1550340 $Y=1576560
X607 5208 5393 5400 1 3 NAND2X2 $T=1626900 1612240 0 0 $X=1626898 $Y=1611838
X608 5933 402 5935 1 3 NAND2X2 $T=1765500 1521520 0 0 $X=1765498 $Y=1521118
X609 6623 6629 6660 1 3 NAND2X2 $T=1949640 1481200 0 180 $X=1946340 $Y=1475760
X610 580 6705 6681 1 3 NAND2X2 $T=1958880 1531600 0 180 $X=1955580 $Y=1526160
X611 6762 584 6740 1 3 NAND2X2 $T=1982640 1561840 1 180 $X=1979340 $Y=1561438
X612 590 6779 6773 1 3 NAND2X2 $T=1987260 1511440 0 180 $X=1983960 $Y=1506000
X613 600 6974 6928 1 3 NAND2X2 $T=2029500 1511440 0 180 $X=2026200 $Y=1506000
X614 601 6944 6941 1 3 NAND2X2 $T=2027520 1491280 0 0 $X=2027518 $Y=1490878
X615 7006 7050 7040 1 3 NAND2X2 $T=2057220 1491280 1 0 $X=2057218 $Y=1485840
X616 7073 7069 7051 1 3 NAND2X2 $T=2061180 1551760 0 180 $X=2057880 $Y=1546320
X617 7824 659 7707 1 3 NAND2X2 $T=2248620 1501360 1 0 $X=2248618 $Y=1495920
X618 7926 663 7864 1 3 NAND2X2 $T=2270400 1491280 1 0 $X=2270398 $Y=1485840
X619 7991 670 671 1 3 NAND2X2 $T=2291520 1430800 0 0 $X=2291518 $Y=1430398
X620 687 8207 8134 1 3 NAND2X2 $T=2348940 1440880 0 0 $X=2348938 $Y=1440478
X621 2420 3 2427 2473 1 2475 AOI21X4 $T=896940 1491280 0 0 $X=896938 $Y=1490878
X622 2622 3 2632 2704 1 2699 AOI21X4 $T=951720 1461040 0 0 $X=951718 $Y=1460638
X623 138 3 2833 2827 1 2743 AOI21X4 $T=991980 1592080 1 180 $X=985380 $Y=1591678
X624 4350 3 343 4347 1 4474 AOI21X4 $T=1380720 1551760 0 0 $X=1380718 $Y=1551358
X625 4812 3 4687 4830 1 373 AOI21X4 $T=1488300 1481200 0 0 $X=1488298 $Y=1480798
X626 5208 3 5399 5462 1 5401 AOI21X4 $T=1642740 1602160 1 0 $X=1642738 $Y=1596720
X627 6683 3 6663 6704 1 6772 AOI21X4 $T=1960200 1491280 1 0 $X=1960198 $Y=1485840
X628 6781 3 6818 6776 1 6878 AOI21X4 $T=1995180 1481200 0 0 $X=1995178 $Y=1480798
X629 6781 3 6818 6776 1 6931 AOI21X4 $T=1996500 1481200 1 0 $X=1996498 $Y=1475760
X630 7359 3 7467 7471 1 7446 AOI21X4 $T=2168760 1481200 0 180 $X=2162160 $Y=1475760
X631 7428 3 7426 7526 1 7511 AOI21X4 $T=2173380 1521520 0 0 $X=2173378 $Y=1521118
X632 7471 3 7528 7587 1 7576 AOI21X4 $T=2188560 1471120 1 0 $X=2188558 $Y=1465680
X633 7655 3 7786 7801 1 656 AOI21X4 $T=2236080 1491280 1 0 $X=2236078 $Y=1485840
X634 7683 3 7874 7879 1 661 AOI21X4 $T=2253240 1450960 1 0 $X=2253238 $Y=1445520
X635 2477 3 2533 1 2550 AND2X2 $T=922680 1450960 1 0 $X=922678 $Y=1445520
X636 2534 3 2515 1 2546 AND2X2 $T=923340 1481200 0 0 $X=923338 $Y=1480798
X637 2724 3 2686 1 2685 AND2X2 $T=953700 1521520 1 180 $X=951060 $Y=1521118
X638 179 3 3157 1 178 AND2X2 $T=1073160 1430800 1 180 $X=1070520 $Y=1430398
X639 197 3 233 1 3588 AND2X2 $T=1178100 1531600 1 0 $X=1178098 $Y=1526160
X640 197 3 265 1 3855 AND2X2 $T=1241460 1440880 1 0 $X=1241458 $Y=1435440
X641 4054 3 4096 1 3955 AND2X2 $T=1309440 1511440 1 180 $X=1306800 $Y=1511038
X642 4414 3 4394 1 4402 AND2X2 $T=1390620 1491280 1 180 $X=1387980 $Y=1490878
X643 355 3 346 1 4597 AND2X2 $T=1437480 1440880 1 0 $X=1437478 $Y=1435440
X644 4594 3 4683 1 4543 AND2X2 $T=1440120 1481200 0 180 $X=1437480 $Y=1475760
X645 4684 3 4683 1 4590 AND2X2 $T=1450680 1471120 1 180 $X=1448040 $Y=1470718
X646 4751 3 4683 1 4693 AND2X2 $T=1469160 1461040 0 180 $X=1466520 $Y=1455600
X647 368 3 4683 1 4817 AND2X2 $T=1479720 1450960 1 0 $X=1479718 $Y=1445520
X648 355 3 363 1 4770 AND2X2 $T=1483680 1430800 1 180 $X=1481040 $Y=1430398
X649 370 3 378 1 4898 AND2X2 $T=1500840 1521520 0 0 $X=1500838 $Y=1521118
X650 392 3 397 1 5151 AND2X2 $T=1564200 1592080 1 180 $X=1561560 $Y=1591678
X651 5201 3 404 1 5127 AND2X2 $T=1571460 1582000 0 180 $X=1568820 $Y=1576560
X652 5298 3 5315 1 5039 AND2X2 $T=1609080 1571920 0 180 $X=1606440 $Y=1566480
X653 5431 3 5421 1 5496 AND2X2 $T=1636800 1501360 1 0 $X=1636798 $Y=1495920
X654 5293 3 421 1 5267 AND2X2 $T=1657260 1440880 0 0 $X=1657258 $Y=1440478
X655 5698 3 192 1 5696 AND2X2 $T=1702800 1491280 0 180 $X=1700160 $Y=1485840
X656 484 3 468 1 6029 AND2X2 $T=1803780 1430800 1 180 $X=1801140 $Y=1430398
X657 484 3 509 1 516 AND2X2 $T=1828860 1430800 0 0 $X=1828858 $Y=1430398
X658 484 3 489 1 6191 AND2X2 $T=1830180 1440880 0 0 $X=1830178 $Y=1440478
X659 6215 3 521 1 6190 AND2X2 $T=1835460 1440880 0 180 $X=1832820 $Y=1435440
X660 544 3 545 1 6362 AND2X2 $T=1895520 1521520 0 0 $X=1895518 $Y=1521118
X661 6584 3 569 1 6357 AND2X2 $T=1941060 1612240 0 0 $X=1941058 $Y=1611838
X662 6683 3 6681 1 6686 AND2X2 $T=1958220 1481200 1 0 $X=1958218 $Y=1475760
X663 584 3 586 1 6754 AND2X2 $T=1981980 1541680 0 180 $X=1979340 $Y=1536240
X664 6773 3 6774 1 6768 AND2X2 $T=1985280 1491280 1 180 $X=1982640 $Y=1490878
X665 7012 3 7006 1 7005 AND2X2 $T=2049960 1491280 0 180 $X=2047320 $Y=1485840
X666 7467 3 7397 1 7363 AND2X2 $T=2148960 1481200 0 180 $X=2146320 $Y=1475760
X667 7813 3 657 1 7866 AND2X2 $T=2252580 1602160 0 0 $X=2252578 $Y=1601758
X668 7861 3 7882 1 7860 AND2X2 $T=2256540 1531600 0 180 $X=2253900 $Y=1526160
X669 8115 3 8134 1 8118 AND2X2 $T=2329800 1440880 1 180 $X=2327160 $Y=1440478
X670 739 3 9080 1 9097 AND2X2 $T=2570040 1602160 1 0 $X=2570038 $Y=1596720
X671 2421 1 111 3 2419 NAND2X4 $T=894960 1521520 1 180 $X=890340 $Y=1521118
X672 4054 1 4061 3 4083 NAND2X4 $T=1300200 1571920 0 0 $X=1300198 $Y=1571518
X673 4489 1 4558 3 356 NAND2X4 $T=1424940 1491280 0 0 $X=1424938 $Y=1490878
X674 4688 1 4686 3 335 NAND2X4 $T=1453320 1592080 1 180 $X=1448700 $Y=1591678
X675 4748 1 4747 3 4721 NAND2X4 $T=1469820 1501360 1 180 $X=1465200 $Y=1500958
X676 4686 1 4780 3 366 NAND2X4 $T=1475100 1602160 1 0 $X=1475098 $Y=1596720
X677 5026 1 388 3 5023 NAND2X4 $T=1542420 1582000 0 180 $X=1537800 $Y=1576560
X678 5129 1 392 3 5026 NAND2X4 $T=1547040 1582000 0 180 $X=1542420 $Y=1576560
X679 5711 1 5534 3 5625 NAND2X4 $T=1707420 1491280 1 0 $X=1707418 $Y=1485840
X680 5176 1 5568 3 472 NAND2X4 $T=1744380 1602160 0 0 $X=1744378 $Y=1601758
X681 581 1 578 3 6629 NAND2X4 $T=1966140 1521520 0 180 $X=1961520 $Y=1516080
X682 6683 1 6623 3 6756 NAND2X4 $T=1968780 1481200 1 0 $X=1968778 $Y=1475760
X683 6739 1 6761 3 6758 NAND2X4 $T=1982640 1551760 1 180 $X=1978020 $Y=1551358
X684 2476 1687 1 3 2533 OR2X2 $T=910800 1450960 1 0 $X=910798 $Y=1445520
X685 1929 2500 1 3 2534 OR2X2 $T=915420 1481200 0 0 $X=915418 $Y=1480798
X686 126 125 1 3 2632 OR2X2 $T=965580 1461040 1 180 $X=962940 $Y=1460638
X687 137 135 1 3 2772 OR2X2 $T=990000 1481200 1 180 $X=987360 $Y=1480798
X688 150 147 1 3 145 OR2X2 $T=1002540 1541680 0 180 $X=999900 $Y=1536240
X689 172 163 1 3 3038 OR2X2 $T=1050720 1481200 1 180 $X=1048080 $Y=1480798
X690 3193 3190 1 3 3157 OR2X2 $T=1085700 1450960 1 180 $X=1083060 $Y=1450558
X691 245 242 1 3 3582 OR2X2 $T=1192620 1592080 1 180 $X=1189980 $Y=1591678
X692 291 242 1 3 3827 OR2X2 $T=1246740 1592080 1 180 $X=1244100 $Y=1591678
X693 302 304 1 3 3834 OR2X2 $T=1279740 1592080 1 180 $X=1277100 $Y=1591678
X694 314 4036 1 3 4101 OR2X2 $T=1302180 1501360 1 0 $X=1302178 $Y=1495920
X695 322 242 1 3 4015 OR2X2 $T=1306800 1612240 0 180 $X=1304160 $Y=1606800
X696 4057 2966 1 3 4131 OR2X2 $T=1310760 1571920 0 0 $X=1310758 $Y=1571518
X697 4097 2213 1 3 4166 OR2X2 $T=1320000 1551760 0 0 $X=1319998 $Y=1551358
X698 330 304 1 3 3585 OR2X2 $T=1322640 1592080 1 180 $X=1320000 $Y=1591678
X699 3037 4146 1 3 4097 OR2X2 $T=1323960 1561840 1 180 $X=1321320 $Y=1561438
X700 85 4101 1 3 4287 OR2X2 $T=1328580 1501360 1 0 $X=1328578 $Y=1495920
X701 329 247 1 3 4014 OR2X2 $T=1331880 1612240 1 180 $X=1329240 $Y=1611838
X702 4041 333 1 3 4248 OR2X2 $T=1345080 1561840 0 0 $X=1345078 $Y=1561438
X703 359 361 1 3 4730 OR2X2 $T=1457280 1551760 0 0 $X=1457278 $Y=1551358
X704 4723 4917 1 3 4835 OR2X2 $T=1508760 1582000 0 180 $X=1506120 $Y=1576560
X705 417 5199 1 3 405 OR2X2 $T=1576740 1430800 1 180 $X=1574100 $Y=1430398
X706 5152 5200 1 3 5195 OR2X2 $T=1605120 1501360 1 0 $X=1605118 $Y=1495920
X707 5326 5220 1 3 5361 OR2X2 $T=1636800 1551760 0 0 $X=1636798 $Y=1551358
X708 449 5646 1 3 5618 OR2X2 $T=1694220 1531600 0 0 $X=1694218 $Y=1531198
X709 5539 5497 1 3 5579 OR2X2 $T=1696860 1450960 1 0 $X=1696858 $Y=1445520
X710 302 537 1 3 6356 OR2X2 $T=1869120 1612240 1 0 $X=1869118 $Y=1606800
X711 537 250 1 3 6435 OR2X2 $T=1895520 1602160 0 0 $X=1895518 $Y=1601758
X712 537 329 1 3 6556 OR2X2 $T=1925880 1612240 1 0 $X=1925878 $Y=1606800
X713 537 330 1 3 6580 OR2X2 $T=1934460 1592080 0 0 $X=1934458 $Y=1591678
X714 537 248 1 3 6584 OR2X2 $T=1934460 1612240 0 0 $X=1934458 $Y=1611838
X715 572 566 1 3 6555 OR2X2 $T=1937760 1602160 0 180 $X=1935120 $Y=1596720
X716 576 6695 1 3 6585 OR2X2 $T=1962180 1582000 1 180 $X=1959540 $Y=1581598
X717 576 577 1 3 6443 OR2X2 $T=1962180 1602160 0 180 $X=1959540 $Y=1596720
X718 590 6779 1 3 6774 OR2X2 $T=1987260 1501360 0 180 $X=1984620 $Y=1495920
X719 554 596 1 3 6942 OR2X2 $T=2021580 1541680 0 0 $X=2021578 $Y=1541278
X720 609 7075 1 3 7073 OR2X2 $T=2065800 1551760 1 0 $X=2065798 $Y=1546320
X721 624 623 1 3 7222 OR2X2 $T=2119260 1582000 1 180 $X=2116620 $Y=1581598
X722 7365 7331 1 3 7307 OR2X2 $T=2134440 1521520 0 180 $X=2131800 $Y=1516080
X723 7444 638 1 3 633 OR2X2 $T=2160840 1612240 1 180 $X=2158200 $Y=1611838
X724 7490 7530 1 3 7445 OR2X2 $T=2180640 1561840 0 180 $X=2178000 $Y=1556400
X725 7555 7557 1 3 7426 OR2X2 $T=2192520 1531600 1 0 $X=2192518 $Y=1526160
X726 7684 7647 1 3 7646 OR2X2 $T=2201760 1592080 1 180 $X=2199120 $Y=1591678
X727 648 7670 1 3 7467 OR2X2 $T=2212320 1450960 1 180 $X=2209680 $Y=1450558
X728 653 7684 1 3 7729 OR2X2 $T=2224860 1592080 1 180 $X=2222220 $Y=1591678
X729 7791 654 1 3 7757 OR2X2 $T=2235420 1592080 0 180 $X=2232780 $Y=1586640
X730 7881 660 1 3 7815 OR2X2 $T=2257860 1582000 1 180 $X=2255220 $Y=1581598
X731 7946 7945 1 3 7861 OR2X2 $T=2277660 1531600 0 180 $X=2275020 $Y=1526160
X732 722 706 1 3 8733 OR2X2 $T=2498100 1491280 1 180 $X=2495460 $Y=1490878
X733 597 720 1 3 8809 OR2X2 $T=2515260 1501360 1 180 $X=2512620 $Y=1500958
X734 9084 9046 1 3 743 OR2X2 $T=2571360 1440880 1 0 $X=2571358 $Y=1435440
X735 9103 9102 1 3 742 OR2X2 $T=2575320 1461040 0 180 $X=2572680 $Y=1455600
X736 9080 722 1 3 9162 OR2X2 $T=2591160 1461040 1 0 $X=2591158 $Y=1455600
X737 9236 9220 1 3 753 OR2X2 $T=2605680 1461040 1 0 $X=2605678 $Y=1455600
X738 27 1 3 34 1569 NAND2XL $T=666600 1511440 1 0 $X=666598 $Y=1506000
X739 1636 1 3 34 1760 NAND2XL $T=711480 1511440 0 0 $X=711478 $Y=1511038
X740 34 1 3 1781 1822 NAND2XL $T=725340 1511440 0 0 $X=725338 $Y=1511038
X741 3177 1 3 3157 3158 NAND2XL $T=1075140 1450960 1 180 $X=1073160 $Y=1450558
X742 4507 1 3 4478 4559 NAND2XL $T=1422300 1511440 1 0 $X=1422298 $Y=1506000
X743 4685 1 3 4598 4603 NAND2XL $T=1442760 1511440 0 180 $X=1440780 $Y=1506000
X744 4779 1 3 4727 4846 NAND2XL $T=1477080 1541680 1 0 $X=1477078 $Y=1536240
X745 5103 1 3 5025 5152 NAND2XL $T=1586640 1501360 0 180 $X=1584660 $Y=1495920
X746 5352 1 3 5298 394 NAND2XL $T=1617660 1561840 1 180 $X=1615680 $Y=1561438
X747 5357 1 3 404 5269 NAND2XL $T=1623600 1501360 0 0 $X=1623598 $Y=1500958
X748 439 1 3 5521 444 NAND2XL $T=1683000 1450960 0 180 $X=1681020 $Y=1445520
X749 5646 1 3 449 5627 NAND2XL $T=1688280 1531600 1 180 $X=1686300 $Y=1531198
X750 5627 1 3 5618 447 NAND2XL $T=1688280 1551760 1 180 $X=1686300 $Y=1551358
X751 439 1 3 5509 5539 NAND2XL $T=1691580 1461040 1 0 $X=1691578 $Y=1455600
X752 5697 1 3 450 5699 NAND2XL $T=1702140 1450960 1 0 $X=1702138 $Y=1445520
X753 591 1 3 6762 6807 NAND2XL $T=1994520 1561840 1 180 $X=1992540 $Y=1561438
X754 567 1 3 571 7120 NAND2XL $T=2083620 1511440 0 180 $X=2081640 $Y=1506000
X755 571 1 3 608 7168 NAND2XL $T=2091540 1501360 1 0 $X=2091538 $Y=1495920
X756 7171 1 3 7222 7236 NAND2XL $T=2106720 1582000 1 180 $X=2104740 $Y=1581598
X757 7488 1 3 7443 7373 NAND2XL $T=2164800 1571920 1 180 $X=2162820 $Y=1571518
X758 7512 1 3 7445 7430 NAND2XL $T=2174700 1561840 1 180 $X=2172720 $Y=1561438
X759 7880 1 3 7815 7709 NAND2XL $T=2255880 1571920 0 180 $X=2253900 $Y=1566480
X760 8122 1 3 8157 8121 NAND2XL $T=2327820 1541680 0 180 $X=2325840 $Y=1536240
X761 8304 1 3 8303 8275 NAND2XL $T=2375340 1511440 1 180 $X=2373360 $Y=1511038
X762 8438 1 3 8422 8428 NAND2XL $T=2410980 1501360 1 0 $X=2410978 $Y=1495920
X763 8478 1 3 8471 702 NAND2XL $T=2419560 1440880 0 180 $X=2417580 $Y=1435440
X764 8471 1 3 8424 8510 NAND2XL $T=2425500 1440880 0 0 $X=2425498 $Y=1440478
X765 8738 1 3 8711 721 NAND2XL $T=2497440 1450960 0 180 $X=2495460 $Y=1445520
X766 592 1 3 598 738 NAND2XL $T=2572680 1612240 1 180 $X=2570700 $Y=1611838
X767 9102 1 3 9103 9117 NAND2XL $T=2573340 1450960 1 0 $X=2573338 $Y=1445520
X768 94 103 1 3 INVX4 $T=873180 1551760 0 0 $X=873178 $Y=1551358
X769 2475 2446 1 3 INVX4 $T=901560 1471120 1 180 $X=898920 $Y=1470718
X770 3627 231 1 3 INVX4 $T=1190640 1551760 0 180 $X=1188000 $Y=1546320
X771 4474 4475 1 3 INVX4 $T=1401180 1541680 0 0 $X=1401178 $Y=1541278
X772 5102 4831 1 3 INVX4 $T=1550340 1592080 1 180 $X=1547700 $Y=1591678
X773 5319 5462 1 3 INVX4 $T=1634820 1592080 0 0 $X=1634818 $Y=1591678
X774 5626 417 1 3 INVX4 $T=1688940 1440880 0 180 $X=1686300 $Y=1435440
X775 5899 5933 1 3 INVX4 $T=1756920 1511440 0 0 $X=1756918 $Y=1511038
X776 5698 5898 1 3 INVX4 $T=1762860 1481200 0 0 $X=1762858 $Y=1480798
X777 5967 476 1 3 INVX4 $T=1772760 1481200 0 0 $X=1772758 $Y=1480798
X778 480 484 1 3 INVX4 $T=1789260 1461040 1 0 $X=1789258 $Y=1455600
X779 554 545 1 3 INVX4 $T=1896840 1551760 1 0 $X=1896838 $Y=1546320
X780 6629 6663 1 3 INVX4 $T=1955580 1491280 0 180 $X=1952940 $Y=1485840
X781 6721 6683 1 3 INVX4 $T=1974060 1501360 0 0 $X=1974058 $Y=1500958
X782 7329 7312 1 3 INVX4 $T=2132460 1561840 0 0 $X=2132458 $Y=1561438
X783 1817 67 3 1823 1765 1 AOI21X1 $T=729300 1582000 0 0 $X=729298 $Y=1581598
X784 2686 2687 3 2688 2623 1 AOI21X1 $T=951720 1511440 0 0 $X=951718 $Y=1511038
X785 2765 2687 3 2762 2758 1 AOI21X1 $T=973500 1511440 0 180 $X=970860 $Y=1506000
X786 2726 2771 3 2773 2782 1 AOI21X1 $T=973500 1561840 1 0 $X=973498 $Y=1556400
X787 99 2905 3 2908 2845 1 AOI21X1 $T=1001880 1571920 1 0 $X=1001878 $Y=1566480
X788 3157 177 3 180 3128 1 AOI21X1 $T=1073160 1450960 0 180 $X=1070520 $Y=1445520
X789 3292 3229 3 3306 3321 1 AOI21X1 $T=1106160 1481200 0 0 $X=1106158 $Y=1480798
X790 194 170 3 3335 3292 1 AOI21X1 $T=1118700 1481200 1 180 $X=1116060 $Y=1480798
X791 4802 4727 3 4795 4803 1 AOI21X1 $T=1483680 1521520 0 0 $X=1483678 $Y=1521118
X792 394 5064 3 5006 5061 1 AOI21X1 $T=1549680 1592080 0 180 $X=1547040 $Y=1586640
X793 5133 396 3 5101 5100 1 AOI21X1 $T=1552980 1511440 1 180 $X=1550340 $Y=1511038
X794 5152 5148 3 5101 5132 1 AOI21X1 $T=1563540 1501360 0 180 $X=1560900 $Y=1495920
X795 387 5256 3 5257 412 1 AOI21X1 $T=1589280 1592080 1 0 $X=1589278 $Y=1586640
X796 5324 5315 3 4744 5257 1 AOI21X1 $T=1602480 1592080 0 180 $X=1599840 $Y=1586640
X797 404 5219 3 5354 5294 1 AOI21X1 $T=1622280 1551760 1 0 $X=1622278 $Y=1546320
X798 429 427 3 5399 432 1 AOI21X1 $T=1626240 1602160 0 0 $X=1626238 $Y=1601758
X799 5430 5513 3 5516 5536 1 AOI21X1 $T=1657920 1582000 1 0 $X=1657918 $Y=1576560
X800 427 5006 3 5698 5543 1 AOI21X1 $T=1716660 1501360 0 0 $X=1716658 $Y=1500958
X801 519 518 3 6193 6187 1 AOI21X1 $T=1835460 1571920 0 180 $X=1832820 $Y=1566480
X802 500 235 3 6292 6291 1 AOI21X1 $T=1856580 1602160 0 180 $X=1853940 $Y=1596720
X803 542 538 3 6362 6325 1 AOI21X1 $T=1873740 1521520 1 180 $X=1871100 $Y=1521118
X804 7006 7038 3 7068 7010 1 AOI21X1 $T=2060520 1501360 1 0 $X=2060518 $Y=1495920
X805 7443 7369 3 7425 7424 1 AOI21X1 $T=2156880 1571920 1 180 $X=2154240 $Y=1571518
X806 7425 7445 3 7474 7449 1 AOI21X1 $T=2165460 1561840 1 0 $X=2165458 $Y=1556400
X807 7815 7732 3 7789 7790 1 AOI21X1 $T=2240700 1582000 0 180 $X=2238060 $Y=1576560
X808 658 7813 3 7795 7811 1 AOI21X1 $T=2245980 1602160 1 180 $X=2243340 $Y=1601758
X809 8062 8064 3 8061 8052 1 AOI21X1 $T=2308680 1511440 0 180 $X=2306040 $Y=1506000
X810 8051 667 3 8067 8086 1 AOI21X1 $T=2306700 1592080 1 0 $X=2306698 $Y=1586640
X811 8065 672 3 8069 8006 1 AOI21X1 $T=2307360 1612240 1 0 $X=2307358 $Y=1606800
X812 8137 8064 3 8154 8166 1 AOI21X1 $T=2331120 1501360 0 0 $X=2331118 $Y=1500958
X813 8154 8200 3 8230 8229 1 AOI21X1 $T=2350920 1511440 1 0 $X=2350918 $Y=1506000
X814 8440 8560 3 8562 709 1 AOI21X1 $T=2444640 1440880 0 0 $X=2444638 $Y=1440478
X815 8786 724 3 8804 725 1 AOI21X1 $T=2504700 1430800 0 0 $X=2504698 $Y=1430398
X816 1780 1565 1 1798 3 1961 OAI21X2 $T=724020 1491280 1 0 $X=724018 $Y=1485840
X817 2419 2394 1 2363 3 2473 OAI21X2 $T=900240 1501360 1 0 $X=900238 $Y=1495920
X818 4726 4800 1 4815 3 4830 OAI21X2 $T=1485660 1481200 1 0 $X=1485658 $Y=1475760
X819 5162 5061 1 5102 3 400 OAI21X2 $T=1564200 1592080 0 180 $X=1558920 $Y=1586640
X820 6928 6946 1 6941 3 7038 OAI21X2 $T=2031480 1481200 1 180 $X=2026200 $Y=1480798
X821 7511 7570 1 7576 3 7683 OAI21X2 $T=2187900 1481200 1 0 $X=2187898 $Y=1475760
X822 7783 7754 1 7766 3 7867 OAI21X2 $T=2243340 1461040 1 0 $X=2243338 $Y=1455600
X823 7707 7794 1 7864 3 7801 OAI21X2 $T=2248620 1491280 1 0 $X=2248618 $Y=1485840
X824 8134 684 1 8186 3 686 OAI21X2 $T=2347620 1440880 1 0 $X=2347618 $Y=1435440
X825 2379 2495 2518 1 3 XNOR2X4 $T=906180 1521520 0 0 $X=906178 $Y=1521118
X826 4241 334 340 1 3 XNOR2X4 $T=1346400 1471120 1 0 $X=1346398 $Y=1465680
X827 6664 6682 579 1 3 XNOR2X4 $T=1955580 1450960 1 0 $X=1955578 $Y=1445520
X828 7040 7039 605 1 3 XNOR2X4 $T=2056560 1461040 0 180 $X=2045340 $Y=1455600
X829 7051 7041 603 1 3 XNOR2X4 $T=2058540 1511440 0 180 $X=2047320 $Y=1506000
X830 8938 8931 7980 1 3 XNOR2X4 $T=2537040 1561840 0 180 $X=2525820 $Y=1556400
X831 1721 1 1669 1654 3 51 OAI21X4 $T=697620 1491280 1 180 $X=690360 $Y=1490878
X832 70 1 1863 1839 3 66 OAI21X4 $T=739860 1571920 0 0 $X=739858 $Y=1571518
X833 2395 1 2496 2419 3 2495 OAI21X4 $T=909480 1531600 0 180 $X=902220 $Y=1526160
X834 2498 1 2475 2509 3 116 OAI21X4 $T=906840 1450960 0 0 $X=906838 $Y=1450558
X835 2723 1 2699 2725 3 123 OAI21X4 $T=957000 1440880 1 0 $X=956998 $Y=1435440
X836 2770 1 2743 2727 3 2622 OAI21X4 $T=968220 1481200 1 180 $X=960960 $Y=1480798
X837 4524 1 344 351 3 4550 OAI21X4 $T=1417680 1592080 1 0 $X=1417678 $Y=1586640
X838 4585 1 4599 4685 3 4687 OAI21X4 $T=1446720 1501360 0 0 $X=1446718 $Y=1500958
X839 4227 1 4745 377 3 375 OAI21X4 $T=1495560 1612240 0 0 $X=1495558 $Y=1611838
X840 5331 1 5354 396 3 358 OAI21X4 $T=1614360 1531600 1 0 $X=1614358 $Y=1526160
X841 5897 1 5898 5534 3 5912 OAI21X4 $T=1754280 1491280 1 0 $X=1754278 $Y=1485840
X842 313 1 5947 5935 3 474 OAI21X4 $T=1770780 1551760 1 180 $X=1763520 $Y=1551358
X843 6666 1 6615 6629 3 6682 OAI21X4 $T=1958880 1471120 0 0 $X=1958878 $Y=1470718
X844 6756 1 6615 6772 3 6760 OAI21X4 $T=1979340 1471120 1 0 $X=1979338 $Y=1465680
X845 6772 1 6787 6773 3 6776 OAI21X4 $T=1989240 1481200 1 180 $X=1981980 $Y=1480798
X846 6930 1 6931 6928 3 6945 OAI21X4 $T=2030160 1471120 1 0 $X=2030158 $Y=1465680
X847 7013 1 6991 7036 3 7039 OAI21X4 $T=2047320 1461040 0 0 $X=2047318 $Y=1460638
X848 626 1 7328 627 3 7329 OAI21X4 $T=2131140 1612240 0 0 $X=2131138 $Y=1611838
X849 7253 1 7429 7449 3 7428 OAI21X4 $T=2154900 1551760 0 0 $X=2154898 $Y=1551358
X850 7668 1 7360 7648 3 7655 OAI21X4 $T=2206380 1511440 0 180 $X=2199120 $Y=1506000
X851 2705 1 47 3 CLKBUFX8 $T=964920 1582000 0 0 $X=964918 $Y=1581598
X852 2708 1 31 3 CLKBUFX8 $T=964920 1612240 0 0 $X=964918 $Y=1611838
X853 3097 1 82 3 CLKBUFX8 $T=1050720 1592080 0 180 $X=1046100 $Y=1586640
X854 3179 1 49 3 CLKBUFX8 $T=1085040 1612240 1 0 $X=1085038 $Y=1606800
X855 3288 1 40 3 CLKBUFX8 $T=1105500 1602160 0 180 $X=1100880 $Y=1596720
X856 3590 1 222 3 CLKBUFX8 $T=1184040 1450960 0 180 $X=1179420 $Y=1445520
X857 3628 1 214 3 CLKBUFX8 $T=1194600 1531600 0 0 $X=1194598 $Y=1531198
X858 232 1 234 3 CLKBUFX8 $T=1199880 1511440 0 0 $X=1199878 $Y=1511038
X859 3841 1 190 3 CLKBUFX8 $T=1241460 1582000 1 180 $X=1236840 $Y=1581598
X860 3922 1 188 3 CLKBUFX8 $T=1259280 1430800 1 180 $X=1254660 $Y=1430398
X861 3969 1 217 3 CLKBUFX8 $T=1277760 1491280 0 180 $X=1273140 $Y=1485840
X862 4139 1 256 3 CLKBUFX8 $T=1321980 1612240 0 180 $X=1317360 $Y=1606800
X863 4135 1 325 3 CLKBUFX8 $T=1327260 1471120 0 0 $X=1327258 $Y=1470718
X864 335 1 4139 3 CLKBUFX8 $T=1348380 1612240 1 0 $X=1348378 $Y=1606800
X865 4369 1 309 3 CLKBUFX8 $T=1378080 1440880 1 0 $X=1378078 $Y=1435440
X866 7287 1 4855 3 CLKBUFX8 $T=2122560 1481200 1 180 $X=2117940 $Y=1480798
X867 1835 1813 3 1 65 XOR2X2 $T=733260 1541680 1 180 $X=726660 $Y=1541278
X868 117 2516 3 1 2740 XOR2X2 $T=913440 1612240 1 0 $X=913438 $Y=1606800
X869 2685 2687 3 1 2444 XOR2X2 $T=955680 1531600 0 180 $X=949080 $Y=1526160
X870 485 563 3 1 574 XOR2X2 $T=1925220 1491280 0 0 $X=1925218 $Y=1490878
X871 6754 6757 3 1 585 XOR2X2 $T=1976040 1531600 1 0 $X=1976038 $Y=1526160
X872 6807 6799 3 1 587 XOR2X2 $T=1994520 1531600 0 180 $X=1987920 $Y=1526160
X873 7363 7359 3 1 7342 XOR2X2 $T=2144340 1481200 1 180 $X=2137740 $Y=1480798
X874 7448 7446 3 1 7423 XOR2X2 $T=2160840 1481200 1 180 $X=2154240 $Y=1480798
X875 7810 7806 3 1 6996 XOR2X2 $T=2245320 1531600 1 180 $X=2238720 $Y=1531198
X876 7860 7856 3 1 6974 XOR2X2 $T=2251920 1521520 1 180 $X=2245320 $Y=1521118
X877 7899 7896 3 1 6944 XOR2X2 $T=2263800 1511440 1 180 $X=2257200 $Y=1511038
X878 8070 8066 3 1 7991 XOR2X2 $T=2310660 1440880 0 180 $X=2304060 $Y=1435440
X879 8118 676 3 1 7926 XOR2X2 $T=2323200 1450960 0 180 $X=2316600 $Y=1445520
X880 104 1 2304 3 INVX2 $T=879120 1561840 1 0 $X=879118 $Y=1556400
X881 2902 1 2938 3 INVX2 $T=1014420 1461040 1 0 $X=1014418 $Y=1455600
X882 169 1 163 3 INVX2 $T=1064580 1501360 0 180 $X=1062600 $Y=1495920
X883 187 1 177 3 INVX2 $T=1086360 1531600 1 180 $X=1084380 $Y=1531198
X884 225 1 211 3 INVX2 $T=1376760 1592080 0 0 $X=1376758 $Y=1591678
X885 289 1 227 3 INVX2 $T=1405140 1602160 0 0 $X=1405138 $Y=1601758
X886 306 1 316 3 INVX2 $T=1431540 1602160 1 0 $X=1431538 $Y=1596720
X887 270 1 255 3 INVX2 $T=1432860 1592080 0 0 $X=1432858 $Y=1591678
X888 240 1 259 3 INVX2 $T=1432860 1612240 0 0 $X=1432858 $Y=1611838
X889 235 1 213 3 INVX2 $T=1443420 1612240 1 0 $X=1443418 $Y=1606800
X890 582 1 6757 3 INVX2 $T=1970760 1541680 1 180 $X=1968780 $Y=1541278
X891 7655 1 7608 3 INVX2 $T=2206380 1491280 0 0 $X=2206378 $Y=1490878
X892 1721 3 1 1801 INVXL $T=727320 1501360 1 0 $X=727318 $Y=1495920
X893 49 3 1 121 INVXL $T=933900 1602160 1 0 $X=933898 $Y=1596720
X894 80 3 1 2728 INVXL $T=966240 1561840 1 180 $X=964920 $Y=1561438
X895 47 3 1 2966 INVXL $T=1019700 1571920 0 0 $X=1019698 $Y=1571518
X896 40 3 1 3551 INVXL $T=1163580 1592080 0 0 $X=1163578 $Y=1591678
X897 231 3 1 3602 INVXL $T=1178100 1481200 0 0 $X=1178098 $Y=1480798
X898 231 3 1 230 INVXL $T=1183380 1430800 1 180 $X=1182060 $Y=1430398
X899 4687 3 1 4725 INVXL $T=1461900 1481200 0 0 $X=1461898 $Y=1480798
X900 378 3 1 4795 INVXL $T=1497540 1521520 1 180 $X=1496220 $Y=1521118
X901 5104 3 1 390 INVXL $T=1533840 1551760 0 180 $X=1532520 $Y=1546320
X902 403 3 1 5162 INVXL $T=1562880 1571920 0 180 $X=1561560 $Y=1566480
X903 5247 3 1 5219 INVXL $T=1595220 1571920 1 0 $X=1595218 $Y=1566480
X904 5315 3 1 425 INVXL $T=1608420 1592080 0 0 $X=1608418 $Y=1591678
X905 5236 3 1 5293 INVXL $T=1660560 1471120 0 0 $X=1660558 $Y=1470718
X906 383 3 1 443 INVXL $T=1668480 1461040 0 0 $X=1668478 $Y=1460638
X907 4745 3 1 5693 INVXL $T=1692240 1582000 0 0 $X=1692238 $Y=1581598
X908 6038 3 1 6028 INVXL $T=1795200 1440880 0 180 $X=1793880 $Y=1435440
X909 529 3 1 503 INVXL $T=1845360 1582000 0 180 $X=1844040 $Y=1576560
X910 531 3 1 525 INVXL $T=1848000 1592080 0 180 $X=1846680 $Y=1586640
X911 8085 3 1 8062 INVXL $T=2310660 1521520 1 180 $X=2309340 $Y=1521118
X912 8089 3 1 8061 INVXL $T=2313300 1521520 0 180 $X=2311980 $Y=1516080
X913 8440 3 1 8427 INVXL $T=2405040 1440880 1 180 $X=2403720 $Y=1440478
X914 8478 3 1 8476 INVXL $T=2418240 1450960 1 180 $X=2416920 $Y=1450558
X915 8497 3 1 8471 INVXL $T=2425500 1450960 0 180 $X=2424180 $Y=1445520
X916 5158 399 407 3 5207 4728 1 AOI31X1 $T=1579380 1592080 0 180 $X=1576080 $Y=1586640
X917 4744 5247 5038 3 5198 5273 1 AOI31X1 $T=1586640 1582000 0 0 $X=1586638 $Y=1581598
X918 5990 490 491 3 487 6034 1 AOI31X1 $T=1793220 1602160 0 0 $X=1793218 $Y=1601758
X919 6116 495 497 3 487 6039 1 AOI31X1 $T=1799820 1582000 1 180 $X=1796520 $Y=1581598
X920 7861 7862 7856 3 7865 7806 1 AOI31X1 $T=2250600 1531600 0 0 $X=2250598 $Y=1531198
X921 1597 1601 3 1 50 XNOR2X2 $T=674520 1511440 1 0 $X=674518 $Y=1506000
X922 1784 1785 3 1 61 XNOR2X2 $T=722040 1450960 0 180 $X=714780 $Y=1445520
X923 2806 2805 3 1 127 XNOR2X2 $T=982080 1612240 1 180 $X=974820 $Y=1611838
X924 528 6509 3 1 612 XNOR2X2 $T=2059200 1430800 0 0 $X=2059198 $Y=1430398
X925 7290 7289 3 1 4617 XNOR2X2 $T=2124540 1521520 1 180 $X=2117280 $Y=1521118
X926 7751 7748 3 1 7287 XNOR2X2 $T=2230140 1491280 0 180 $X=2222880 $Y=1485840
X927 7875 7867 3 1 7824 XNOR2X2 $T=2256540 1461040 1 180 $X=2249280 $Y=1460638
X928 1742 1740 1 3 1723 XOR2X1 $T=711480 1592080 1 180 $X=706200 $Y=1591678
X929 1767 1765 1 3 1661 XOR2X1 $T=715440 1551760 0 180 $X=710160 $Y=1546320
X930 2624 2623 1 3 2421 XOR2X1 $T=945780 1521520 1 180 $X=940500 $Y=1521118
X931 2700 2699 1 3 2476 XOR2X1 $T=956340 1440880 1 180 $X=951060 $Y=1440478
X932 2759 2758 1 3 2347 XOR2X1 $T=972180 1501360 1 180 $X=966900 $Y=1500958
X933 3031 168 1 3 164 XOR2X1 $T=1042800 1471120 1 180 $X=1037520 $Y=1470718
X934 3127 3128 1 3 173 XOR2X1 $T=1064580 1450960 0 180 $X=1059300 $Y=1445520
X935 3225 183 1 3 3193 XOR2X1 $T=1094940 1440880 1 180 $X=1089660 $Y=1440478
X936 186 188 1 3 3225 XOR2X1 $T=1102860 1440880 0 180 $X=1097580 $Y=1435440
X937 4395 344 1 3 3415 XOR2X1 $T=1387980 1592080 0 180 $X=1382700 $Y=1586640
X938 4404 4417 1 3 4487 XOR2X1 $T=1390620 1561840 0 0 $X=1390618 $Y=1561438
X939 347 348 1 3 4490 XOR2X1 $T=1401180 1612240 0 0 $X=1401178 $Y=1611838
X940 4544 4509 1 3 3425 XOR2X1 $T=1422300 1551760 1 180 $X=1417020 $Y=1551358
X941 4603 4599 1 3 4594 XOR2X1 $T=1442760 1501360 0 180 $X=1437480 $Y=1495920
X942 4720 4725 1 3 4684 XOR2X1 $T=1463880 1481200 0 180 $X=1458600 $Y=1475760
X943 364 4730 1 3 362 XOR2X1 $T=1469160 1551760 1 180 $X=1463880 $Y=1551358
X944 4795 4792 1 3 367 XOR2X1 $T=1482360 1521520 0 180 $X=1477080 $Y=1516080
X945 6600 571 1 3 5646 XOR2X1 $T=1945020 1521520 1 180 $X=1939740 $Y=1521118
X946 7311 7312 1 3 7293 XOR2X1 $T=2131140 1561840 0 180 $X=2125860 $Y=1556400
X947 7430 7424 1 3 634 XOR2X1 $T=2157540 1582000 0 180 $X=2152260 $Y=1576560
X948 640 7472 1 3 7490 XOR2X1 $T=2164800 1440880 0 0 $X=2164798 $Y=1440478
X949 7529 7360 1 3 7269 XOR2X1 $T=2180640 1511440 1 180 $X=2175360 $Y=1511038
X950 7549 642 1 3 7531 XOR2X1 $T=2185920 1440880 1 180 $X=2180640 $Y=1440478
X951 7756 7754 1 3 7712 XOR2X1 $T=2230800 1461040 1 180 $X=2225520 $Y=1460638
X952 8053 8052 1 3 7933 XOR2X1 $T=2306040 1501360 1 180 $X=2300760 $Y=1500958
X953 8167 8166 1 3 7960 XOR2X1 $T=2339040 1481200 1 180 $X=2333760 $Y=1480798
X954 8292 695 1 3 8235 XOR2X1 $T=2374020 1461040 0 180 $X=2368740 $Y=1455600
X955 8734 8731 1 3 7881 XOR2X1 $T=2496780 1582000 1 180 $X=2491500 $Y=1581598
X956 594 575 1 3 8734 XOR2X1 $T=2504700 1582000 1 180 $X=2499420 $Y=1581598
X957 9105 9086 1 3 7946 XOR2X1 $T=2575320 1541680 0 180 $X=2570040 $Y=1536240
X958 9129 597 1 3 9086 XOR2X1 $T=2583240 1561840 1 180 $X=2577960 $Y=1561438
X959 9129 592 1 3 746 XOR2X1 $T=2580600 1612240 0 0 $X=2580598 $Y=1611838
X960 1560 3 7 1562 1 NOR2BX1 $T=669240 1471120 1 180 $X=666600 $Y=1470718
X961 63 3 62 1740 1 NOR2BX1 $T=718080 1612240 0 180 $X=715440 $Y=1606800
X962 1875 3 1849 1835 1 NOR2BX1 $T=739200 1551760 1 180 $X=736560 $Y=1551358
X963 4779 3 371 4802 1 NOR2BX1 $T=1488960 1541680 0 0 $X=1488958 $Y=1541278
X964 5038 3 5050 5051 1 NOR2BX1 $T=1549020 1551760 1 180 $X=1546380 $Y=1551358
X965 8882 3 8857 730 1 NOR2BX1 $T=2523180 1430800 1 180 $X=2520540 $Y=1430398
X966 575 3 711 9171 1 NOR2BX1 $T=2597760 1551760 1 180 $X=2595120 $Y=1551358
X967 31 36 1587 45 3 1 1598 ADDFX2 $T=663960 1561840 1 0 $X=663958 $Y=1556400
X968 49 32 40 1564 3 1 22 ADDFX2 $T=679140 1592080 0 180 $X=665280 $Y=1586640
X969 1583 47 1564 1581 3 1 35 ADDFX2 $T=681780 1571920 1 180 $X=667920 $Y=1571518
X970 2124 2016 2001 1993 3 1 1930 ADDFX2 $T=784740 1561840 1 180 $X=770880 $Y=1561438
X971 2085 2049 2028 74 3 1 1927 ADDFX2 $T=791340 1461040 0 180 $X=777480 $Y=1455600
X972 2062 2050 2029 1997 3 1 1856 ADDFX2 $T=791340 1481200 1 180 $X=777480 $Y=1480798
X973 2182 2126 2086 1960 3 1 75 ADDFX2 $T=807180 1602160 0 180 $X=793320 $Y=1596720
X974 82 81 80 78 3 1 2084 ADDFX2 $T=811140 1450960 0 180 $X=797280 $Y=1445520
X975 2169 2084 2123 79 3 1 77 ADDFX2 $T=811800 1430800 1 180 $X=797940 $Y=1430398
X976 2129 2138 2125 2123 3 1 2085 ADDFX2 $T=811800 1471120 1 180 $X=797940 $Y=1470718
X977 85 82 81 2069 3 1 2122 ADDFX2 $T=812460 1531600 1 180 $X=798600 $Y=1531198
X978 2122 2142 2130 2051 3 1 2001 ADDFX2 $T=813780 1541680 1 180 $X=799920 $Y=1541278
X979 2127 2155 2128 2028 3 1 2029 ADDFX2 $T=816420 1481200 1 180 $X=802560 $Y=1480798
X980 92 87 83 2129 3 1 2127 ADDFX2 $T=816420 1491280 1 180 $X=802560 $Y=1490878
X981 80 81 84 2049 3 1 2128 ADDFX2 $T=817080 1461040 0 180 $X=803220 $Y=1455600
X982 2139 89 2141 1928 3 1 1959 ADDFX2 $T=817080 1592080 0 180 $X=803220 $Y=1586640
X983 82 85 88 2167 3 1 2126 ADDFX2 $T=803880 1561840 1 0 $X=803878 $Y=1556400
X984 98 2159 86 2139 3 1 2086 ADDFX2 $T=819060 1612240 1 180 $X=805200 $Y=1611838
X985 2187 2167 2158 2124 3 1 2141 ADDFX2 $T=822360 1561840 1 180 $X=808500 $Y=1561438
X986 2209 2196 2184 91 3 1 2169 ADDFX2 $T=832260 1450960 0 180 $X=818400 $Y=1445520
X987 2199 2185 2194 2062 3 1 2030 ADDFX2 $T=835560 1511440 1 180 $X=821700 $Y=1511038
X988 104 92 93 2185 3 1 2130 ADDFX2 $T=835560 1531600 0 180 $X=821700 $Y=1526160
X989 97 101 94 2184 3 1 2125 ADDFX2 $T=836220 1471120 1 180 $X=822360 $Y=1470718
X990 100 101 97 2016 3 1 2187 ADDFX2 $T=839520 1592080 0 180 $X=825660 $Y=1586640
X991 94 97 90 2155 3 1 2194 ADDFX2 $T=840840 1491280 1 180 $X=826980 $Y=1490878
X992 2211 102 2208 2182 3 1 95 ADDFX2 $T=840840 1602160 0 180 $X=826980 $Y=1596720
X993 106 105 102 2050 3 1 2199 ADDFX2 $T=842820 1521520 0 180 $X=828960 $Y=1516080
X994 105 106 2213 2142 3 1 2158 ADDFX2 $T=844140 1561840 0 180 $X=830280 $Y=1556400
X995 81 85 2304 2208 3 1 109 ADDFX2 $T=864600 1602160 1 180 $X=850740 $Y=1601758
X996 568 612 628 630 3 1 635 ADDFX2 $T=2127840 1430800 0 0 $X=2127838 $Y=1430398
X997 682 679 8130 8119 3 1 7990 ADDFX2 $T=2335740 1582000 1 180 $X=2321880 $Y=1581598
X998 677 678 680 8155 3 1 8130 ADDFX2 $T=2322540 1592080 0 0 $X=2322538 $Y=1591678
X999 8155 681 8131 8122 3 1 8101 ADDFX2 $T=2336400 1561840 1 180 $X=2322540 $Y=1561438
X1000 8236 577 689 8196 3 1 8131 ADDFX2 $T=2360160 1561840 0 180 $X=2346300 $Y=1556400
X1001 8196 690 8242 8247 3 1 8157 ADDFX2 $T=2348940 1551760 0 0 $X=2348938 $Y=1551358
X1002 688 8231 8243 8248 3 1 8242 ADDFX2 $T=2348940 1582000 1 0 $X=2348938 $Y=1576560
X1003 678 691 6661 8249 3 1 8243 ADDFX2 $T=2348940 1602160 1 0 $X=2348938 $Y=1596720
X1004 8248 8249 696 8304 3 1 8245 ADDFX2 $T=2370060 1561840 1 0 $X=2370058 $Y=1556400
X1005 699 8349 8355 8345 3 1 8303 ADDFX2 $T=2399760 1541680 1 180 $X=2385900 $Y=1541278
X1006 693 8374 588 8349 3 1 697 ADDFX2 $T=2400420 1602160 1 180 $X=2386560 $Y=1601758
X1007 8368 8381 8425 8438 3 1 8353 ADDFX2 $T=2393820 1521520 0 0 $X=2393818 $Y=1521118
X1008 698 592 566 8381 3 1 8442 ADDFX2 $T=2393820 1571920 1 0 $X=2393818 $Y=1566480
X1009 8442 700 8382 8368 3 1 8355 ADDFX2 $T=2407680 1571920 1 180 $X=2393820 $Y=1571518
X1010 712 678 703 8469 3 1 8382 ADDFX2 $T=2428140 1592080 1 180 $X=2414280 $Y=1591678
X1011 8477 8489 8509 8511 3 1 8422 ADDFX2 $T=2418900 1521520 0 0 $X=2418898 $Y=1521118
X1012 8487 8469 8495 8477 3 1 8425 ADDFX2 $T=2433420 1551760 0 180 $X=2419560 $Y=1546320
X1013 705 598 6695 8489 3 1 8487 ADDFX2 $T=2433420 1571920 0 180 $X=2419560 $Y=1566480
X1014 710 693 677 8530 3 1 8495 ADDFX2 $T=2447280 1582000 1 180 $X=2433420 $Y=1581598
X1015 706 698 577 8615 3 1 8563 ADDFX2 $T=2440680 1541680 1 0 $X=2440678 $Y=1536240
X1016 8616 8615 8552 8551 3 1 8508 ADDFX2 $T=2455200 1501360 1 180 $X=2441340 $Y=1500958
X1017 8625 8530 8563 8552 3 1 8509 ADDFX2 $T=2455200 1531600 0 180 $X=2441340 $Y=1526160
X1018 712 594 711 8626 3 1 8625 ADDFX2 $T=2471040 1571920 1 180 $X=2457180 $Y=1571518
X1019 8626 8644 8653 8654 3 1 8616 ADDFX2 $T=2458500 1561840 0 0 $X=2458498 $Y=1561438
X1020 8684 8683 8654 8671 3 1 8627 ADDFX2 $T=2484900 1511440 1 180 $X=2471040 $Y=1511038
X1021 8681 8700 8714 8711 3 1 8682 ADDFX2 $T=2478960 1481200 1 0 $X=2478958 $Y=1475760
X1022 8729 8699 8701 8681 3 1 8684 ADDFX2 $T=2493480 1531600 1 180 $X=2479620 $Y=1531198
X1023 705 720 717 8701 3 1 8653 ADDFX2 $T=2496120 1571920 1 180 $X=2482260 $Y=1571518
X1024 8728 8733 8740 8785 3 1 8714 ADDFX2 $T=2492820 1481200 0 0 $X=2492818 $Y=1480798
X1025 727 712 8780 8740 3 1 8683 ADDFX2 $T=2510640 1511440 1 180 $X=2496780 $Y=1511038
X1026 8859 8805 8785 8781 3 1 8738 ADDFX2 $T=2513940 1471120 1 180 $X=2500080 $Y=1470718
X1027 723 722 727 8831 3 1 8848 ADDFX2 $T=2504040 1521520 0 0 $X=2504038 $Y=1521118
X1028 8832 710 566 8805 3 1 8700 ADDFX2 $T=2517900 1551760 0 180 $X=2504040 $Y=1546320
X1029 8809 706 8848 8853 3 1 8859 ADDFX2 $T=2508000 1491280 0 0 $X=2507998 $Y=1490878
X1030 726 720 8831 8858 3 1 8899 ADDFX2 $T=2508660 1531600 1 0 $X=2508658 $Y=1526160
X1031 8853 8879 8899 8910 3 1 8883 ADDFX2 $T=2518560 1481200 0 0 $X=2518558 $Y=1480798
X1032 8992 8907 8858 732 3 1 8884 ADDFX2 $T=2537700 1471120 1 180 $X=2523840 $Y=1470718
X1033 592 597 8832 8907 3 1 8879 ADDFX2 $T=2541000 1521520 0 180 $X=2527140 $Y=1516080
X1034 8832 592 8780 8976 3 1 9045 ADDFX2 $T=2539680 1531600 0 0 $X=2539678 $Y=1531198
X1035 8976 677 9043 9046 3 1 737 ADDFX2 $T=2542320 1511440 1 0 $X=2542318 $Y=1506000
X1036 9045 9042 9008 736 3 1 735 ADDFX2 $T=2559480 1450960 0 180 $X=2545620 $Y=1445520
X1037 711 723 9004 9008 3 1 8992 ADDFX2 $T=2560800 1481200 0 180 $X=2546940 $Y=1475760
X1038 723 722 9080 9107 3 1 9110 ADDFX2 $T=2564100 1491280 0 0 $X=2564098 $Y=1490878
X1039 9080 715 598 9078 3 1 9043 ADDFX2 $T=2580600 1501360 1 180 $X=2566740 $Y=1500958
X1040 9078 577 9110 9102 3 1 9084 ADDFX2 $T=2568060 1481200 0 0 $X=2568058 $Y=1480798
X1041 711 715 9162 747 3 1 748 ADDFX2 $T=2583240 1450960 1 0 $X=2583238 $Y=1445520
X1042 9107 717 9176 9220 3 1 9103 ADDFX2 $T=2588520 1491280 0 0 $X=2588518 $Y=1490878
X1043 9170 598 9219 751 3 1 9236 ADDFX2 $T=2595120 1461040 0 0 $X=2595118 $Y=1460638
X1044 72 1945 1 3 73 XNOR2X1 $T=757680 1511440 0 0 $X=757678 $Y=1511038
X1045 1770 1739 1 3 76 XNOR2X1 $T=789360 1511440 0 0 $X=789358 $Y=1511038
X1046 83 99 1 3 2209 XNOR2X1 $T=841500 1450960 0 180 $X=836220 $Y=1445520
X1047 102 108 1 3 2138 XNOR2X1 $T=850740 1471120 1 180 $X=845460 $Y=1470718
X1048 2621 2622 1 3 2500 XNOR2X1 $T=945780 1481200 0 180 $X=940500 $Y=1475760
X1049 2832 136 1 3 133 XNOR2X1 $T=990660 1471120 0 180 $X=985380 $Y=1465680
X1050 4351 4354 1 3 4532 XNOR2X1 $T=1372140 1551760 1 0 $X=1372138 $Y=1546320
X1051 4402 4437 1 3 4510 XNOR2X1 $T=1398540 1491280 1 0 $X=1398538 $Y=1485840
X1052 4508 4491 1 3 3521 XNOR2X1 $T=1411740 1551760 1 180 $X=1406460 $Y=1551358
X1053 4559 4475 1 3 4583 XNOR2X1 $T=1427580 1511440 1 0 $X=1427578 $Y=1506000
X1054 361 4727 1 3 360 XNOR2X1 $T=1463880 1531600 0 180 $X=1458600 $Y=1526160
X1055 4801 4799 1 3 4751 XNOR2X1 $T=1485000 1461040 1 180 $X=1479720 $Y=1460638
X1056 4851 4846 1 3 372 XNOR2X1 $T=1498200 1531600 1 180 $X=1492920 $Y=1531198
X1057 451 452 1 3 456 XNOR2X1 $T=1694220 1551760 1 0 $X=1694218 $Y=1546320
X1058 7109 7108 1 3 610 XNOR2X1 $T=2078340 1521520 1 180 $X=2073060 $Y=1521118
X1059 607 608 1 3 7139 XNOR2X1 $T=2080980 1471120 0 0 $X=2080978 $Y=1470718
X1060 7131 7133 1 3 615 XNOR2X1 $T=2083620 1450960 1 0 $X=2083618 $Y=1445520
X1061 7236 618 1 3 619 XNOR2X1 $T=2104740 1602160 0 0 $X=2104738 $Y=1601758
X1062 622 621 1 3 620 XNOR2X1 $T=2117940 1430800 1 180 $X=2112660 $Y=1430398
X1063 629 7342 1 3 7311 XNOR2X1 $T=2141700 1541680 1 180 $X=2136420 $Y=1541278
X1064 7373 7369 1 3 625 XNOR2X1 $T=2146320 1571920 1 180 $X=2141040 $Y=1571518
X1065 7427 7428 1 3 7444 XNOR2X1 $T=2154900 1541680 1 0 $X=2154898 $Y=1536240
X1066 646 645 1 3 7555 XNOR2X1 $T=2191200 1430800 1 180 $X=2185920 $Y=1430398
X1067 7958 7957 1 3 7671 XNOR2X1 $T=2282280 1612240 1 180 $X=2277000 $Y=1611838
X1068 8087 8064 1 3 8063 XNOR2X1 $T=2313960 1501360 1 180 $X=2308680 $Y=1500958
X1069 8262 8259 1 3 8088 XNOR2X1 $T=2364780 1481200 1 180 $X=2359500 $Y=1480798
X1070 8357 8326 1 3 8334 XNOR2X1 $T=2392500 1471120 0 180 $X=2387220 $Y=1465680
X1071 706 722 1 3 8729 XNOR2X1 $T=2498100 1531600 0 180 $X=2492820 $Y=1526160
X1072 720 597 1 3 8728 XNOR2X1 $T=2503380 1501360 1 180 $X=2498100 $Y=1500958
X1073 594 711 1 3 8938 XNOR2X1 $T=2541660 1582000 1 180 $X=2536380 $Y=1581598
X1074 8938 8832 1 3 733 XNOR2X1 $T=2539020 1592080 0 0 $X=2539018 $Y=1591678
X1075 9095 9080 1 3 9105 XNOR2X1 $T=2571360 1551760 1 0 $X=2571358 $Y=1546320
X1076 715 726 1 3 9129 XNOR2X1 $T=2575320 1602160 1 0 $X=2575318 $Y=1596720
X1077 722 9080 1 3 9170 XNOR2X1 $T=2585880 1471120 0 0 $X=2585878 $Y=1470718
X1078 72 130 1 130 3 2986 3021 3037 OAI221XL $T=1045440 1561840 0 180 $X=1040820 $Y=1556400
X1079 242 251 1 248 3 247 3613 3220 OAI221XL $T=1201860 1612240 1 180 $X=1197240 $Y=1611838
X1080 274 276 1 277 3 278 3812 3811 OAI221XL $T=1229580 1481200 0 0 $X=1229578 $Y=1480798
X1081 242 323 1 321 3 247 319 3936 OAI221XL $T=1305480 1612240 1 180 $X=1300860 $Y=1611838
X1082 5025 5251 1 5259 3 5218 5269 5225 OAI221XL $T=1589940 1501360 0 0 $X=1589938 $Y=1500958
X1083 4041 5198 1 398 3 5274 5412 5430 OAI221XL $T=1631520 1582000 1 0 $X=1631518 $Y=1576560
X1084 5236 440 1 5535 3 5539 5544 5448 OAI221XL $T=1660560 1461040 0 0 $X=1660558 $Y=1460638
X1085 5579 436 1 5497 3 444 445 5356 OAI221XL $T=1673760 1440880 1 0 $X=1673758 $Y=1435440
X1086 6326 6325 1 533 3 6207 6245 6307 OAI221XL $T=1863180 1521520 1 180 $X=1858560 $Y=1521118
X1087 39 1583 41 3 1 1587 ADDHXL $T=666600 1571920 1 0 $X=666598 $Y=1566480
X1088 101 2211 100 3 1 2159 ADDHXL $T=836880 1612240 0 180 $X=829620 $Y=1606800
X1089 468 6215 489 3 1 532 ADDHXL $T=1840740 1440880 1 0 $X=1840738 $Y=1435440
X1090 693 8236 692 3 1 8231 ADDHXL $T=2359500 1592080 0 180 $X=2352240 $Y=1586640
X1091 727 9004 598 3 1 9042 ADDHXL $T=2544300 1491280 0 0 $X=2544298 $Y=1490878
X1092 3 1770 56 1781 1 NOR2XL $T=716100 1521520 1 0 $X=716098 $Y=1516080
X1093 3 147 149 2918 1 NOR2XL $T=1006500 1481200 1 0 $X=1006498 $Y=1475760
X1094 3 3038 170 2904 1 NOR2XL $T=1050060 1481200 0 180 $X=1048080 $Y=1475760
X1095 3 5025 313 5046 1 NOR2XL $T=1543740 1511440 0 0 $X=1543738 $Y=1511038
X1096 3 5198 5162 397 1 NOR2XL $T=1568160 1592080 0 180 $X=1566180 $Y=1586640
X1097 3 5113 5152 5357 1 NOR2XL $T=1608420 1491280 0 0 $X=1608418 $Y=1490878
X1098 3 5195 5180 5327 1 NOR2XL $T=1608420 1521520 1 0 $X=1608418 $Y=1516080
X1099 3 401 427 5330 1 NOR2XL $T=1608420 1602160 1 0 $X=1608418 $Y=1596720
X1100 3 409 434 5220 1 NOR2XL $T=1645380 1561840 0 180 $X=1643400 $Y=1556400
X1101 3 436 4531 438 1 NOR2XL $T=1647360 1440880 1 0 $X=1647358 $Y=1435440
X1102 3 5509 442 5521 1 NOR2XL $T=1668480 1450960 0 0 $X=1668478 $Y=1450558
X1103 3 5509 439 5523 1 NOR2XL $T=1688940 1471120 1 0 $X=1688938 $Y=1465680
X1104 3 664 665 8059 1 NOR2XL $T=2296140 1561840 1 0 $X=2296138 $Y=1556400
X1105 3 8780 575 9079 1 NOR2XL $T=2552220 1582000 1 0 $X=2552218 $Y=1576560
X1106 3 575 597 9187 1 NOR2XL $T=2596440 1571920 1 0 $X=2596438 $Y=1566480
X1107 7139 568 7169 1 3 616 XOR3X2 $T=2104740 1471120 1 180 $X=2092860 $Y=1470718
X1108 673 7990 7982 1 3 7652 XOR3X2 $T=2299440 1571920 1 180 $X=2287560 $Y=1571518
X1109 715 756 755 1 3 7791 XOR3X2 $T=2620200 1602160 1 180 $X=2608320 $Y=1601758
X1110 1636 52 3 1651 1 1659 AOI21XL $T=689700 1511440 0 0 $X=689698 $Y=1511038
X1111 4478 4475 3 4477 1 4437 AOI21XL $T=1406460 1511440 0 180 $X=1403820 $Y=1506000
X1112 4227 398 3 399 1 401 AOI21XL $T=1562220 1612240 0 0 $X=1562218 $Y=1611838
X1113 5198 5218 3 4041 1 5130 AOI21XL $T=1578720 1582000 1 180 $X=1576080 $Y=1581598
X1114 5162 419 3 5298 1 5268 AOI21XL $T=1598520 1561840 1 0 $X=1598518 $Y=1556400
X1115 5025 5253 3 5271 1 5329 AOI21XL $T=1607760 1521520 0 0 $X=1607758 $Y=1521118
X1116 5195 5153 3 416 1 5331 AOI21XL $T=1607760 1531600 1 0 $X=1607758 $Y=1526160
X1117 5523 436 3 454 1 5746 AOI21XL $T=1702140 1471120 1 0 $X=1702138 $Y=1465680
X1118 8440 8471 3 8476 1 8486 AOI21XL $T=2417580 1440880 0 0 $X=2417578 $Y=1440478
X1119 1803 66 1814 1 1785 3 OAI2BB1X1 $T=727320 1440880 0 0 $X=727318 $Y=1440478
X1120 72 130 2809 1 2773 3 OAI2BB1X1 $T=980760 1561840 0 0 $X=980758 $Y=1561438
X1121 3226 3424 3321 1 3479 3 OAI2BB1X1 $T=1142460 1461040 1 0 $X=1142458 $Y=1455600
X1122 448 5618 5627 1 451 3 OAI2BB1X1 $T=1686960 1551760 1 0 $X=1686958 $Y=1546320
X1123 6160 6117 6161 1 6210 3 OAI2BB1X1 $T=1822920 1521520 1 0 $X=1822918 $Y=1516080
X1124 577 715 9188 1 749 3 OAI2BB1X1 $T=2597100 1602160 1 0 $X=2597098 $Y=1596720
X1125 1782 1 41 3 1834 NAND2BXL $T=728640 1521520 0 0 $X=728638 $Y=1521118
X1126 1872 1 1862 3 1784 NAND2BXL $T=741840 1450960 0 180 $X=739200 $Y=1445520
X1127 82 1 118 3 2569 NAND2BXL $T=922680 1582000 0 0 $X=922678 $Y=1581598
X1128 108 1 47 3 2936 NAND2BXL $T=1006500 1561840 1 0 $X=1006498 $Y=1556400
X1129 147 1 195 3 3477 NAND2BXL $T=1149060 1430800 0 0 $X=1149058 $Y=1430398
X1130 283 1 281 3 3812 NAND2BXL $T=1240140 1481200 0 0 $X=1240138 $Y=1480798
X1131 4524 1 351 3 4395 NAND2BXL $T=1413060 1592080 0 180 $X=1410420 $Y=1586640
X1132 488 1 486 3 6016 NAND2BXL $T=1793220 1501360 0 0 $X=1793218 $Y=1500958
X1133 528 1 523 3 6245 NAND2BXL $T=1851300 1521520 0 0 $X=1851298 $Y=1521118
X1134 684 1 8186 3 8070 NAND2BXL $T=2343000 1440880 0 180 $X=2340360 $Y=1435440
X1135 58 60 1 3 CLKBUFX3 $T=702900 1471120 0 0 $X=702898 $Y=1470718
X1136 335 338 1 3 CLKBUFX3 $T=1385340 1592080 0 0 $X=1385338 $Y=1591678
X1137 4745 450 1 3 CLKBUFX3 $T=1690260 1582000 1 0 $X=1690258 $Y=1576560
X1138 561 568 1 3 CLKBUFX3 $T=1931820 1511440 1 0 $X=1931818 $Y=1506000
X1139 2689 224 235 237 3 1 3624 AOI2BB2X1 $T=1181400 1612240 1 0 $X=1181398 $Y=1606800
X1140 331 4041 4096 325 3 1 4152 AOI2BB2X1 $T=1330560 1521520 0 180 $X=1325940 $Y=1516080
X1141 506 510 306 500 3 1 6173 AOI2BB2X1 $T=1817640 1602160 1 0 $X=1817638 $Y=1596720
X1142 520 510 500 225 3 1 6188 AOI2BB2X1 $T=1834140 1602160 0 180 $X=1829520 $Y=1596720
X1143 525 510 500 270 3 1 6209 AOI2BB2X1 $T=1842060 1592080 1 180 $X=1837440 $Y=1591678
X1144 514 510 240 500 3 1 6288 AOI2BB2X1 $T=1846020 1602160 1 0 $X=1846018 $Y=1596720
X1145 2069 2051 2030 1878 3 1 1992 ADDFHX1 $T=796620 1521520 1 180 $X=781440 $Y=1521118
X1146 3557 1 3582 3 3585 3230 NAND3X1 $T=1179420 1592080 0 0 $X=1179418 $Y=1591678
X1147 3777 1 3827 3 3834 3342 NAND3X1 $T=1236840 1592080 0 0 $X=1236838 $Y=1591678
X1148 3876 1 4015 3 4014 308 NAND3X1 $T=1288980 1612240 0 0 $X=1288978 $Y=1611838
X1149 5218 1 5274 3 5315 5380 NAND3X1 $T=1614360 1571920 0 0 $X=1614358 $Y=1571518
X1150 407 1 434 3 399 5274 NAND3X1 $T=1638120 1561840 1 180 $X=1635480 $Y=1561438
X1151 6291 1 6435 3 6443 6411 NAND3X1 $T=1895520 1592080 0 0 $X=1895518 $Y=1591678
X1152 542 1 545 3 6498 6541 NAND3X1 $T=1910040 1511440 1 0 $X=1910038 $Y=1506000
X1153 6124 1 6555 3 6556 6538 NAND3X1 $T=1925880 1602160 1 0 $X=1925878 $Y=1596720
X1154 6188 1 6580 3 6585 6665 NAND3X1 $T=1935780 1582000 0 0 $X=1935778 $Y=1581598
X1155 592 597 715 9219 1 3 9176 CMPR32X1 $T=2587200 1511440 0 0 $X=2587198 $Y=1511038
X1156 7646 7686 7685 1 7693 3 AOI2BB1X2 $T=2209680 1592080 1 0 $X=2209678 $Y=1586640
X1157 5274 5038 1 3 5240 OR2X1 $T=1589280 1602160 0 180 $X=1586640 $Y=1596720
X1158 96 3 90 1 CLKINVX3 $T=830280 1450960 0 0 $X=830278 $Y=1450558
X1159 82 3 107 1 CLKINVX3 $T=838860 1571920 0 0 $X=838858 $Y=1571518
X1160 108 3 2213 1 CLKINVX3 $T=863940 1551760 0 0 $X=863938 $Y=1551358
X1161 2743 3 2687 1 CLKINVX3 $T=967560 1521520 0 0 $X=967558 $Y=1521118
X1162 2970 3 3018 1 CLKINVX3 $T=1035540 1491280 1 0 $X=1035538 $Y=1485840
X1163 176 3 110 1 CLKINVX3 $T=1063260 1612240 0 180 $X=1061280 $Y=1606800
X1164 4831 3 4686 1 CLKINVX3 $T=1484340 1592080 1 180 $X=1482360 $Y=1591678
X1165 5115 3 5101 1 CLKINVX3 $T=1555620 1501360 0 180 $X=1553640 $Y=1495920
X1166 5148 3 5164 1 CLKINVX3 $T=1566180 1501360 1 0 $X=1566178 $Y=1495920
X1167 483 3 485 1 CLKINVX3 $T=1785960 1551760 0 0 $X=1785958 $Y=1551358
X1168 6666 3 6623 1 CLKINVX3 $T=1955580 1481200 0 180 $X=1953600 $Y=1475760
X1169 6681 3 6704 1 CLKINVX3 $T=1958220 1491280 1 180 $X=1956240 $Y=1490878
X1170 7012 3 7013 1 CLKINVX3 $T=2049960 1471120 0 0 $X=2049958 $Y=1470718
X1171 7038 3 7036 1 CLKINVX3 $T=2052600 1481200 0 0 $X=2052598 $Y=1480798
X1172 6798 3 566 1 CLKINVX3 $T=2060520 1582000 0 180 $X=2058540 $Y=1576560
X1173 7397 3 7471 1 CLKINVX3 $T=2172720 1471120 0 0 $X=2172718 $Y=1470718
X1174 7671 3 7530 1 CLKINVX3 $T=2195820 1592080 0 180 $X=2193840 $Y=1586640
X1175 652 3 7736 1 CLKINVX3 $T=2220240 1612240 1 0 $X=2220238 $Y=1606800
X1176 658 3 653 1 CLKINVX3 $T=2247960 1612240 1 180 $X=2245980 $Y=1611838
X1177 8278 3 695 1 CLKINVX3 $T=2369400 1481200 0 0 $X=2369398 $Y=1480798
X1178 594 3 588 1 CLKINVX3 $T=2459820 1592080 0 180 $X=2457840 $Y=1586640
X1179 677 3 723 1 CLKINVX3 $T=2502060 1602160 0 180 $X=2500080 $Y=1596720
X1180 566 3 715 1 CLKINVX3 $T=2614920 1592080 0 0 $X=2614918 $Y=1591678
X1181 739 740 3 1 8731 AND2X1 $T=2572680 1592080 0 180 $X=2570040 $Y=1586640
X1182 5220 5158 3 5129 5201 406 1 AOI22X1 $T=1578060 1571920 1 180 $X=1574760 $Y=1571518
X1183 5180 5022 3 413 414 5104 1 AOI22X1 $T=1584000 1531600 1 0 $X=1583998 $Y=1526160
X1184 7109 7119 3 571 567 7153 1 AOI22X1 $T=2087580 1511440 1 0 $X=2087578 $Y=1506000
X1185 461 5734 5525 5734 1 3 5735 OAI2BB2X1 $T=1717320 1521520 1 180 $X=1712700 $Y=1521118
X1186 462 5734 5746 5734 1 3 5773 OAI2BB2X1 $T=1717980 1471120 1 0 $X=1717978 $Y=1465680
X1187 465 5734 5567 5734 1 3 5777 OAI2BB2X1 $T=1719300 1531600 0 0 $X=1719298 $Y=1531198
X1188 370 4803 1 3 369 XNOR2XL $T=1486320 1511440 0 180 $X=1481040 $Y=1506000
X1189 664 665 1 3 7945 XNOR2XL $T=2275020 1561840 1 0 $X=2275018 $Y=1556400
X1190 710 715 1 3 8644 XNOR2XL $T=2486880 1561840 1 180 $X=2481600 $Y=1561438
X1191 597 575 1 3 9270 XNOR2XL $T=2596440 1582000 1 0 $X=2596438 $Y=1576560
X1192 113 2444 112 3 1 OR2X4 $T=898920 1602160 0 180 $X=894960 $Y=1596720
X1193 106 4287 4241 3 1 OR2X4 $T=1349700 1491280 1 0 $X=1349698 $Y=1485840
X1194 355 313 4204 3 1 OR2X4 $T=1432200 1521520 0 180 $X=1428240 $Y=1516080
X1195 4860 4041 4841 3 1 OR2X4 $T=1497540 1582000 1 180 $X=1493580 $Y=1581598
X1196 476 5933 480 3 1 OR2X4 $T=1783320 1461040 0 0 $X=1783318 $Y=1460638
X1197 484 313 487 3 1 OR2X4 $T=1788600 1561840 0 0 $X=1788598 $Y=1561438
X1198 563 483 564 3 1 OR2X4 $T=1927200 1440880 0 0 $X=1927198 $Y=1440478
X1199 582 6740 6739 3 1 OR2X4 $T=1978020 1551760 1 180 $X=1974060 $Y=1551358
X1200 604 6996 7006 3 1 OR2X4 $T=2044680 1531600 1 0 $X=2044678 $Y=1526160
X1201 528 6509 606 3 1 OR2X4 $T=2047980 1430800 0 0 $X=2047978 $Y=1430398
X1202 647 7649 7528 3 1 OR2X4 $T=2203740 1461040 1 180 $X=2199780 $Y=1460638
X1203 7980 7974 7862 3 1 OR2X4 $T=2287560 1541680 1 180 $X=2283600 $Y=1541278
X1204 326 4101 4143 1 3 324 OAI2BB1X4 $T=1324620 1491280 1 180 $X=1318020 $Y=1490878
X1205 6900 7005 7010 1 3 7041 OAI2BB1X4 $T=2045340 1501360 1 0 $X=2045338 $Y=1495920
X1206 651 7866 7811 1 3 7856 OAI2BB1X4 $T=2251920 1602160 1 0 $X=2251918 $Y=1596720
X1207 58 1565 1 3 INVX8 $T=705540 1471120 0 0 $X=705538 $Y=1470718
X1208 4083 198 1 3 INVX8 $T=1305480 1571920 0 0 $X=1305478 $Y=1571518
X1209 389 5006 1 3 INVX8 $T=1529220 1571920 0 0 $X=1529218 $Y=1571518
X1210 6758 6615 1 3 INVX8 $T=1978020 1481200 1 0 $X=1978018 $Y=1475760
X1211 597 711 1 3 INVX8 $T=2594460 1531600 0 0 $X=2594458 $Y=1531198
X1212 4056 314 4040 320 3 1 MX2X4 $T=1298220 1461040 0 0 $X=1298218 $Y=1460638
X1213 7651 7650 7608 4785 3 1 MX2X4 $T=2203080 1501360 0 180 $X=2196480 $Y=1495920
X1214 410 5267 5241 1 5294 5299 3 OAI2BB2X4 $T=1591260 1551760 1 0 $X=1591258 $Y=1546320
X1215 2395 2419 2472 1 3 NAND2BX2 $T=902220 1541680 1 0 $X=902218 $Y=1536240
X1216 4936 5006 4748 1 3 NAND2BX2 $T=1532520 1501360 0 0 $X=1532518 $Y=1500958
X1217 5352 5895 5909 1 3 NAND2BX2 $T=1754280 1571920 0 0 $X=1754278 $Y=1571518
X1218 5912 5899 470 1 3 NAND2BX2 $T=1758240 1531600 1 180 $X=1754280 $Y=1531198
X1219 5913 5006 5899 1 3 NAND2BX2 $T=1758900 1511440 0 180 $X=1754940 $Y=1506000
X1220 6930 6928 6912 1 3 NAND2BX2 $T=2022900 1461040 1 180 $X=2018940 $Y=1460638
X1221 156 157 2954 2902 3 1 OAI2BB1X2 $T=1021680 1450960 0 180 $X=1017060 $Y=1445520
X1222 5038 5071 395 393 3 1 OAI2BB1X2 $T=1552320 1602160 1 180 $X=1547700 $Y=1601758
X1223 5775 427 5176 5895 3 1 OAI2BB1X2 $T=1744380 1571920 0 0 $X=1744378 $Y=1571518
X1224 443 5579 5582 1 3 5734 AND3X1 $T=1674420 1461040 0 0 $X=1674418 $Y=1460638
X1225 2903 136 2904 1 3 142 AND3X2 $T=997260 1471120 1 180 $X=993960 $Y=1470718
X1226 5420 5517 5407 1 3 5537 AND3X2 $T=1658580 1612240 1 0 $X=1658578 $Y=1606800
X1227 7862 7861 7878 1 3 7859 AND3X2 $T=2259180 1541680 1 180 $X=2255880 $Y=1541278
X1228 536 8059 1 3 7974 XOR2XL $T=2311320 1561840 0 180 $X=2306040 $Y=1556400
X1229 3 3604 244 2304 110 1 NAND3X2 $T=1186680 1571920 0 0 $X=1186678 $Y=1571518
X1230 129 128 82 2749 122 3 1 2705 SDFFRHQXL $T=972840 1602160 0 180 $X=956340 $Y=1596720
X1231 129 128 165 167 122 3 1 3097 SDFFRHQXL $T=1036860 1612240 0 0 $X=1036858 $Y=1611838
X1232 129 128 194 3338 122 3 1 3307 SDFFRHQXL $T=1123980 1511440 0 180 $X=1107480 $Y=1506000
X1233 129 128 94 3320 122 3 1 3362 SDFFRHQXL $T=1108140 1561840 0 0 $X=1108138 $Y=1561438
X1234 129 128 96 3340 122 3 1 3234 SDFFRHQXL $T=1124640 1551760 1 180 $X=1108140 $Y=1551358
X1235 129 128 193 3355 122 3 1 3304 SDFFRHQXL $T=1127280 1582000 0 180 $X=1110780 $Y=1576560
X1236 129 128 184 3356 122 3 1 3421 SDFFRHQXL $T=1120020 1501360 1 0 $X=1120018 $Y=1495920
X1237 129 128 195 3391 122 3 1 3344 SDFFRHQXL $T=1137180 1440880 1 180 $X=1120680 $Y=1440478
X1238 129 241 3602 3603 232 3 1 3566 SDFFRHQXL $T=1193280 1501360 0 180 $X=1176780 $Y=1495920
X1239 129 241 201 3520 234 3 1 3548 SDFFRHQXL $T=1195920 1511440 0 180 $X=1179420 $Y=1506000
X1240 129 241 222 246 234 3 1 3598 SDFFRHQXL $T=1202520 1491280 0 180 $X=1186020 $Y=1485840
X1241 129 241 204 249 234 3 1 3601 SDFFRHQXL $T=1205160 1471120 0 180 $X=1188660 $Y=1465680
X1242 129 241 203 252 234 3 1 3590 SDFFRHQXL $T=1207140 1450960 1 180 $X=1190640 $Y=1450558
X1243 129 241 185 3698 232 3 1 3628 SDFFRHQXL $T=1213080 1521520 1 180 $X=1196580 $Y=1521118
X1244 129 241 80 261 232 3 1 3627 SDFFRHQXL $T=1217040 1551760 0 180 $X=1200540 $Y=1546320
X1245 129 241 216 3497 234 3 1 3743 SDFFRHQXL $T=1203180 1501360 0 0 $X=1203178 $Y=1500958
X1246 129 128 281 3837 182 3 1 3906 SDFFRHQXL $T=1235520 1561840 0 0 $X=1235518 $Y=1561438
X1247 129 241 284 3840 232 3 1 3907 SDFFRHQXL $T=1236180 1531600 0 0 $X=1236178 $Y=1531198
X1248 129 128 108 298 182 3 1 3841 SDFFRHQXL $T=1265880 1582000 1 180 $X=1249380 $Y=1581598
X1249 129 128 190 3936 232 3 1 3838 SDFFRHQXL $T=1265880 1612240 1 180 $X=1249380 $Y=1611838
X1250 129 128 303 301 122 3 1 3922 SDFFRHQXL $T=1282380 1430800 1 180 $X=1265880 $Y=1430398
X1251 129 241 188 3965 234 3 1 3969 SDFFRHQXL $T=1267860 1501360 1 0 $X=1267858 $Y=1495920
X1252 129 241 217 3924 234 3 1 294 SDFFRHQXL $T=1269180 1481200 1 0 $X=1269178 $Y=1475760
X1253 129 128 296 3882 122 3 1 285 SDFFRHQXL $T=1290960 1430800 0 0 $X=1290958 $Y=1430398
X1254 129 241 309 4017 122 3 1 296 SDFFRHQXL $T=1290960 1450960 1 0 $X=1290958 $Y=1445520
X1255 332 241 294 4175 234 3 1 4135 SDFFRHQXL $T=1334520 1461040 1 180 $X=1318020 $Y=1460638
X1256 129 241 325 4134 234 3 1 292 SDFFRHQXL $T=1318680 1450960 1 0 $X=1318678 $Y=1445520
X1257 332 241 292 4238 234 3 1 4324 SDFFRHQXL $T=1347060 1450960 1 0 $X=1347058 $Y=1445520
X1258 332 241 346 4319 234 3 1 4369 SDFFRHQXL $T=1393260 1450960 0 180 $X=1376760 $Y=1445520
X1259 332 241 349 4528 234 3 1 346 SDFFRHQXL $T=1422960 1450960 0 180 $X=1406460 $Y=1445520
X1260 332 241 4531 4529 234 3 1 349 SDFFRHQXL $T=1422960 1450960 1 180 $X=1406460 $Y=1450558
X1261 332 241 339 4691 234 3 1 363 SDFFRHQXL $T=1450020 1440880 1 0 $X=1450018 $Y=1435440
X1262 332 241 363 4854 234 3 1 384 SDFFRHQXL $T=1493580 1440880 1 0 $X=1493578 $Y=1435440
X1263 332 241 384 5107 234 3 1 5025 SDFFRHQXL $T=1557600 1440880 1 180 $X=1541100 $Y=1440478
X1264 332 241 5025 5045 234 3 1 5063 SDFFRHQXL $T=1541760 1461040 1 0 $X=1541758 $Y=1455600
X1265 332 241 5113 5323 234 3 1 5103 SDFFRHQXL $T=1603800 1461040 1 0 $X=1603798 $Y=1455600
X1266 428 241 5103 5356 234 3 1 423 SDFFRHQXL $T=1620960 1440880 0 180 $X=1604460 $Y=1435440
X1267 332 241 436 5448 234 3 1 4531 SDFFRHQXL $T=1648680 1461040 0 180 $X=1632180 $Y=1455600
X1268 332 241 5509 5600 234 3 1 436 SDFFRHQXL $T=1682340 1511440 1 0 $X=1682338 $Y=1506000
X1269 332 241 455 5576 234 3 1 5509 SDFFRHQXL $T=1699500 1511440 1 180 $X=1683000 $Y=1511038
X1270 332 464 462 5735 463 3 1 5789 SDFFRHQXL $T=1717320 1511440 0 0 $X=1717318 $Y=1511038
X1271 332 464 461 5777 463 3 1 5747 SDFFRHQXL $T=1733820 1541680 1 180 $X=1717320 $Y=1541278
X1272 332 464 459 5700 463 3 1 5725 SDFFRHQXL $T=1734480 1561840 1 180 $X=1717980 $Y=1561438
X1273 332 464 467 5756 463 3 1 5749 SDFFRHQXL $T=1735140 1602160 1 180 $X=1718640 $Y=1601758
X1274 332 464 453 5773 463 3 1 5812 SDFFRHQXL $T=1722600 1461040 1 0 $X=1722598 $Y=1455600
X1275 332 464 468 5699 463 3 1 5930 SDFFRHQXL $T=1747680 1450960 1 0 $X=1747678 $Y=1445520
X1276 332 464 489 6028 463 3 1 468 SDFFRHQXL $T=1797840 1440880 1 180 $X=1781340 $Y=1440478
X1277 332 464 509 6139 463 3 1 489 SDFFRHQXL $T=1822260 1440880 0 180 $X=1805760 $Y=1435440
X1278 332 464 531 6330 541 3 1 6377 SDFFRHQXL $T=1859880 1571920 1 0 $X=1859878 $Y=1566480
X1279 332 547 6157 6411 541 3 1 6478 SDFFRHQXL $T=1884300 1571920 1 0 $X=1884298 $Y=1566480
X1280 332 464 529 6442 541 3 1 6495 SDFFRHQXL $T=1892880 1561840 1 0 $X=1892878 $Y=1556400
X1281 332 464 575 6665 541 3 1 553 SDFFRHQXL $T=1959540 1551760 1 180 $X=1943040 $Y=1551358
X1282 332 547 592 6801 541 3 1 6881 SDFFRHQXL $T=1992540 1612240 1 0 $X=1992538 $Y=1606800
X1283 332 547 6798 6759 541 3 1 6882 SDFFRHQXL $T=1993200 1592080 1 0 $X=1993198 $Y=1586640
X1284 332 547 597 6808 541 3 1 7070 SDFFRHQXL $T=2018940 1582000 0 0 $X=2018938 $Y=1581598
X1285 1565 3 38 1 BUFX3 $T=667920 1461040 1 0 $X=667918 $Y=1455600
X1286 104 3 87 1 BUFX3 $T=835560 1531600 1 0 $X=835558 $Y=1526160
X1287 36 3 3130 1 BUFX3 $T=1045440 1541680 0 0 $X=1045438 $Y=1541278
X1288 130 3 193 1 BUFX3 $T=1090320 1521520 0 0 $X=1090318 $Y=1521118
X1289 3307 3 184 1 BUFX3 $T=1108800 1501360 1 0 $X=1108798 $Y=1495920
X1290 3362 3 99 1 BUFX3 $T=1126620 1561840 1 0 $X=1126618 $Y=1556400
X1291 3344 3 194 1 BUFX3 $T=1127280 1430800 0 0 $X=1127278 $Y=1430398
X1292 3421 3 201 1 BUFX3 $T=1143120 1501360 0 0 $X=1143118 $Y=1500958
X1293 99 3 218 1 BUFX3 $T=1153020 1541680 0 0 $X=1153018 $Y=1541278
X1294 3548 3 185 1 BUFX3 $T=1171500 1511440 0 180 $X=1168860 $Y=1506000
X1295 3566 3 204 1 BUFX3 $T=1176780 1471120 1 180 $X=1174140 $Y=1470718
X1296 3743 3 192 1 BUFX3 $T=1211760 1481200 1 180 $X=1209120 $Y=1480798
X1297 3906 3 272 1 BUFX3 $T=1242780 1561840 0 180 $X=1240140 $Y=1556400
X1298 3883 3 3881 1 BUFX3 $T=1250700 1511440 1 180 $X=1248060 $Y=1511038
X1299 3907 3 281 1 BUFX3 $T=1259280 1531600 0 0 $X=1259278 $Y=1531198
X1300 128 3 241 1 BUFX3 $T=1265880 1531600 0 0 $X=1265878 $Y=1531198
X1301 5500 3 402 1 BUFX3 $T=1654620 1521520 0 180 $X=1651980 $Y=1516080
X1302 4745 3 446 1 BUFX3 $T=1680360 1602160 0 0 $X=1680358 $Y=1601758
X1303 5725 3 455 1 BUFX3 $T=1710720 1561840 1 180 $X=1708080 $Y=1561438
X1304 5747 3 465 1 BUFX3 $T=1721280 1551760 0 0 $X=1721278 $Y=1551358
X1305 5749 3 459 1 BUFX3 $T=1721280 1602160 1 0 $X=1721278 $Y=1596720
X1306 5789 3 461 1 BUFX3 $T=1726560 1521520 1 180 $X=1723920 $Y=1521118
X1307 5812 3 462 1 BUFX3 $T=1734480 1471120 0 180 $X=1731840 $Y=1465680
X1308 5930 3 453 1 BUFX3 $T=1757580 1440880 0 180 $X=1754940 $Y=1435440
X1309 6377 3 534 1 BUFX3 $T=1873080 1582000 0 180 $X=1870440 $Y=1576560
X1310 6478 3 558 1 BUFX3 $T=1906740 1571920 1 0 $X=1906738 $Y=1566480
X1311 5895 3 560 1 BUFX3 $T=1916640 1582000 0 0 $X=1916638 $Y=1581598
X1312 6882 3 575 1 BUFX3 $T=2000460 1571920 1 180 $X=1997820 $Y=1571518
X1313 6881 3 598 1 BUFX3 $T=2020920 1612240 1 0 $X=2020918 $Y=1606800
X1314 6931 3 6991 1 BUFX3 $T=2031480 1461040 0 0 $X=2031478 $Y=1460638
X1315 7070 3 594 1 BUFX3 $T=2065800 1582000 1 0 $X=2065798 $Y=1576560
X1316 7293 3 4488 1 BUFX3 $T=2110020 1561840 0 180 $X=2107380 $Y=1556400
X1317 7269 3 4637 1 BUFX3 $T=2117940 1511440 1 180 $X=2115300 $Y=1511038
X1318 575 3 722 1 BUFX3 $T=2505360 1541680 1 0 $X=2505358 $Y=1536240
X1319 594 3 9080 1 BUFX3 $T=2554860 1602160 0 0 $X=2554858 $Y=1601758
X1320 285 199 207 3 183 1 3855 3857 AOI221X1 $T=1246740 1430800 1 180 $X=1242120 $Y=1430398
X1321 387 386 385 3 4096 1 328 4936 AOI221X1 $T=1518660 1501360 1 180 $X=1514040 $Y=1500958
X1322 5256 427 5219 3 5326 1 403 5412 AOI221X1 $T=1620960 1582000 1 0 $X=1620958 $Y=1576560
X1323 5521 439 5150 3 402 1 5510 5525 AOI221X1 $T=1662540 1521520 0 180 $X=1657920 $Y=1516080
X1324 5946 414 5945 3 427 1 5465 5913 AOI221X1 $T=1768140 1501360 1 180 $X=1763520 $Y=1500958
X1325 156 221 3477 3 147 3435 1 3437 AOI32XL $T=1152360 1440880 0 180 $X=1147740 $Y=1435440
X1326 3772 267 266 3 262 265 1 3729 AOI32XL $T=1222980 1440880 0 180 $X=1218360 $Y=1435440
X1327 277 278 3812 3 283 282 1 3752 AOI32XL $T=1242780 1481200 0 180 $X=1238160 $Y=1475760
X1328 6085 6121 483 3 6048 494 1 6086 AOI32XL $T=1809060 1521520 1 180 $X=1804440 $Y=1521118
X1329 533 6207 6245 3 528 6231 1 6204 AOI32XL $T=1848000 1521520 1 180 $X=1843380 $Y=1521118
X1330 6289 6230 524 3 6302 501 1 6306 AOI32XL $T=1853940 1461040 0 0 $X=1853938 $Y=1460638
X1331 6361 6355 6157 3 6346 536 1 6304 AOI32XL $T=1872420 1481200 0 180 $X=1867800 $Y=1475760
X1332 1770 32 3 1 CLKINVX4 $T=737220 1531600 0 0 $X=737218 $Y=1531198
X1333 268 271 3 1 CLKINVX4 $T=1224960 1602160 1 0 $X=1224958 $Y=1596720
X1334 4054 4086 3 1 CLKINVX4 $T=1304820 1561840 0 0 $X=1304818 $Y=1561438
X1335 4868 4860 3 1 CLKINVX4 $T=1500180 1582000 0 180 $X=1497540 $Y=1576560
X1336 5726 5711 3 1 CLKINVX4 $T=1711380 1501360 0 180 $X=1708740 $Y=1495920
X1337 5912 5947 3 1 CLKINVX4 $T=1768140 1541680 0 0 $X=1768138 $Y=1541278
X1338 589 6762 3 1 CLKINVX4 $T=1979340 1582000 1 180 $X=1976700 $Y=1581598
X1339 169 197 3 199 185 207 214 3433 1 AOI222X2 $T=1155000 1521520 0 180 $X=1145760 $Y=1516080
X1340 4728 4723 1 4745 4744 3 4749 OAI22X1 $T=1469160 1602160 0 180 $X=1465200 $Y=1596720
X1341 416 5237 1 415 5274 3 5226 OAI22X1 $T=1592580 1612240 1 0 $X=1592578 $Y=1606800
X1342 5512 5535 1 5498 5524 3 5576 OAI22X1 $T=1664520 1501360 0 180 $X=1660560 $Y=1495920
X1343 6162 6187 1 6162 6163 3 6161 OAI22X1 $T=1826880 1561840 0 180 $X=1822920 $Y=1556400
X1344 566 560 1 573 329 3 6658 OAI22X1 $T=1950960 1592080 0 180 $X=1947000 $Y=1586640
X1345 6661 560 1 573 302 3 6801 OAI22X1 $T=1974720 1612240 0 180 $X=1970760 $Y=1606800
X1346 6695 560 1 573 330 3 6759 OAI22X1 $T=1976040 1592080 0 180 $X=1972080 $Y=1586640
X1347 588 560 1 573 307 3 6808 OAI22X1 $T=1983960 1592080 0 180 $X=1980000 $Y=1586640
X1348 1593 3 43 1597 1 NOR2BXL $T=677160 1521520 0 0 $X=677158 $Y=1521118
X1349 82 3 118 2619 1 NOR2BXL $T=939180 1582000 0 0 $X=939178 $Y=1581598
X1350 108 3 47 2908 1 NOR2BXL $T=1013760 1571920 0 180 $X=1011120 $Y=1566480
X1351 184 3 175 3228 1 NOR2BXL $T=1097580 1491280 1 180 $X=1094940 $Y=1490878
X1352 192 3 136 3335 1 NOR2BXL $T=1126620 1481200 1 180 $X=1123980 $Y=1480798
X1353 511 3 512 6175 1 NOR2BXL $T=1822260 1551760 0 0 $X=1822258 $Y=1551358
X1354 475 3 531 6193 1 NOR2BXL $T=1848660 1571920 0 180 $X=1846020 $Y=1566480
X1355 3226 3 3474 3531 1 3533 NOR3BX1 $T=1163580 1450960 0 0 $X=1163578 $Y=1450558
X1356 6160 3 6099 6120 1 6205 NOR3BX1 $T=1822920 1511440 1 0 $X=1822918 $Y=1506000
X1357 185 3 163 3231 1 3228 3226 AOI211X1 $T=1096920 1481200 0 180 $X=1093620 $Y=1475760
X1358 3796 3 3799 3764 1 3811 3774 AOI211X1 $T=1230900 1461040 1 0 $X=1230898 $Y=1455600
X1359 5129 3 391 5130 1 5134 4917 AOI211X1 $T=1558920 1582000 1 0 $X=1558918 $Y=1576560
X1360 5149 3 396 5046 1 5101 5147 AOI211X1 $T=1564860 1511440 1 180 $X=1561560 $Y=1511038
X1361 5237 3 398 411 1 409 408 AOI211X1 $T=1582020 1602160 1 180 $X=1578720 $Y=1601758
X1362 5200 3 5253 5197 1 5149 5251 AOI211X1 $T=1591260 1511440 1 180 $X=1587960 $Y=1511038
X1363 5494 3 5523 5521 1 396 5512 AOI211X1 $T=1661880 1491280 0 180 $X=1658580 $Y=1485840
X1364 402 3 5254 438 1 5521 5567 AOI211X1 $T=1666500 1521520 1 0 $X=1666498 $Y=1516080
X1365 515 3 514 6178 1 6175 6160 AOI211X1 $T=1831500 1551760 1 180 $X=1828200 $Y=1551358
X1366 6324 3 6322 6206 1 6307 6286 AOI211X1 $T=1861200 1511440 0 180 $X=1857900 $Y=1506000
X1367 8938 3 8990 8993 1 711 8901 AOI211X1 $T=2544960 1551760 0 0 $X=2544958 $Y=1551358
X1368 3018 163 2973 1 169 3052 3 3008 OAI32X1 $T=1042800 1501360 1 0 $X=1042798 $Y=1495920
X1369 3228 185 163 1 184 172 3 3229 OAI32X1 $T=1097580 1491280 0 180 $X=1092960 $Y=1485840
X1370 3335 194 170 1 192 191 3 3306 OAI32X1 $T=1119360 1491280 0 180 $X=1114740 $Y=1485840
X1371 3774 3748 3479 1 3533 3479 3 264 OAI32X1 $T=1221660 1461040 0 180 $X=1217040 $Y=1455600
X1372 5194 5352 5153 1 5298 419 3 5354 OAI32X1 $T=1613040 1541680 0 0 $X=1613038 $Y=1541278
X1373 6175 515 514 1 511 517 3 6163 OAI32X1 $T=1830180 1561840 1 0 $X=1830178 $Y=1556400
X1374 6286 6216 6210 1 6205 6210 3 6214 OAI32X1 $T=1841400 1511440 0 180 $X=1836780 $Y=1506000
X1375 6193 519 518 1 475 525 3 6162 OAI32X1 $T=1837440 1571920 0 0 $X=1837438 $Y=1571518
X1376 6362 538 542 1 544 545 3 6326 OAI32X1 $T=1880340 1521520 0 0 $X=1880338 $Y=1521118
X1377 44 1569 1 3 48 1601 AOI2BB1X1 $T=676500 1501360 0 0 $X=676498 $Y=1500958
X1378 72 2986 1 3 2782 3021 AOI2BB1X1 $T=1026960 1561840 1 0 $X=1026958 $Y=1556400
X1379 404 5207 1 3 411 435 AOI2BB1X1 $T=1636140 1602160 0 0 $X=1636138 $Y=1601758
X1380 307 537 1 3 6542 6494 AOI2BB1X1 $T=1924560 1592080 1 180 $X=1921260 $Y=1591678
X1381 7736 7735 1 3 7732 7727 AOI2BB1X1 $T=2224860 1582000 0 180 $X=2221560 $Y=1576560
X1382 9187 566 1 3 9171 8993 AOI2BB1X1 $T=2597760 1561840 0 180 $X=2594460 $Y=1556400
X1383 207 204 3 199 194 197 3399 168 1 AOI222X1 $T=1142460 1471120 1 180 $X=1137180 $Y=1470718
X1384 39 198 3 200 104 3415 3390 206 1 AOI222X1 $T=1138500 1561840 0 0 $X=1138498 $Y=1561438
X1385 200 82 3 209 206 3413 3395 118 1 AOI222X1 $T=1144440 1582000 1 180 $X=1139160 $Y=1581598
X1386 199 201 3 203 207 197 3408 159 1 AOI222X1 $T=1139820 1481200 0 0 $X=1139818 $Y=1480798
X1387 31 198 3 200 94 3425 3397 206 1 AOI222X1 $T=1139820 1551760 0 0 $X=1139818 $Y=1551358
X1388 49 198 3 200 105 210 3429 206 1 AOI222X1 $T=1139820 1612240 1 0 $X=1139818 $Y=1606800
X1389 197 175 3 199 184 207 3434 216 1 AOI222X1 $T=1142460 1491280 0 0 $X=1142458 $Y=1490878
X1390 207 217 3 199 192 136 3480 197 1 AOI222X1 $T=1155000 1481200 1 180 $X=1149720 $Y=1480798
X1391 206 3521 3 80 200 3514 3492 40 1 AOI222X1 $T=1164240 1551760 1 180 $X=1158960 $Y=1551358
X1392 197 269 3 199 272 273 3792 207 1 AOI222X1 $T=1223640 1531600 1 0 $X=1223638 $Y=1526160
X1393 199 281 3 190 207 197 3845 283 1 AOI222X1 $T=1237500 1521520 0 0 $X=1237498 $Y=1521118
X1394 197 277 3 199 294 295 3919 207 1 AOI222X1 $T=1252680 1481200 1 0 $X=1252678 $Y=1475760
X1395 287 197 3 199 296 188 3986 207 1 AOI222X1 $T=1255980 1450960 1 0 $X=1255978 $Y=1445520
X1396 197 288 3 199 292 207 3937 297 1 AOI222X1 $T=1257300 1450960 0 0 $X=1257298 $Y=1450558
X1397 153 149 2902 1 3 143 XNOR3X2 $T=1009800 1450960 1 180 $X=997920 $Y=1450558
X1398 7153 608 571 1 3 611 XNOR3X2 $T=2089560 1541680 1 180 $X=2077680 $Y=1541278
X1399 288 3 3877 287 286 3799 1 AOI22XL $T=1246080 1450960 1 180 $X=1242780 $Y=1450558
X1400 32 3 4061 4112 96 4288 1 AOI22XL $T=1313400 1521520 0 0 $X=1313398 $Y=1521118
X1401 41 3 4061 4112 193 4224 1 AOI22XL $T=1313400 1531600 0 0 $X=1313398 $Y=1531198
X1402 3130 3 4061 4112 218 4120 1 AOI22XL $T=1313400 1541680 0 0 $X=1313398 $Y=1541278
X1403 5180 3 402 396 5149 5131 1 AOI22XL $T=1564860 1521520 0 180 $X=1561560 $Y=1516080
X1404 5129 3 5219 5220 328 5071 1 AOI22XL $T=1579380 1561840 1 180 $X=1576080 $Y=1561438
X1405 5256 3 427 403 5326 5390 1 AOI22XL $T=1621620 1592080 1 0 $X=1621618 $Y=1586640
X1406 5327 3 5419 5361 414 5431 1 AOI22XL $T=1632180 1511440 0 0 $X=1632178 $Y=1511038
X1407 5246 3 5521 5577 5318 5582 1 AOI22XL $T=1671780 1471120 0 0 $X=1671778 $Y=1470718
X1408 557 3 6381 539 6364 6322 1 AOI22XL $T=1884300 1501360 1 180 $X=1881000 $Y=1500958
X1409 163 2973 1 175 3 3041 AOI2BB1XL $T=1065240 1491280 1 180 $X=1061940 $Y=1490878
X1410 286 287 1 292 3 3877 AOI2BB1XL $T=1254000 1450960 1 180 $X=1250700 $Y=1450558
X1411 5152 5218 1 328 3 5227 AOI2BB1XL $T=1584660 1501360 1 180 $X=1581360 $Y=1500958
X1412 6364 539 1 540 3 6381 AOI2BB1XL $T=1873080 1501360 0 0 $X=1873078 $Y=1500958
X1413 9086 9095 1 9080 3 9082 AOI2BB1XL $T=2575980 1551760 0 0 $X=2575978 $Y=1551358
X1414 172 3018 3 3031 1 3041 166 AOI211X2 $T=1046760 1491280 0 180 $X=1040820 $Y=1485840
X1415 3234 94 1 3 BUFX4 $T=1096260 1551760 1 180 $X=1092960 $Y=1551358
X1416 3304 96 1 3 BUFX4 $T=1108800 1541680 1 180 $X=1105500 $Y=1541278
X1417 3601 203 1 3 BUFX4 $T=1191960 1461040 1 0 $X=1191958 $Y=1455600
X1418 3598 216 1 3 BUFX4 $T=1195920 1491280 0 0 $X=1195918 $Y=1490878
X1419 4324 339 1 3 BUFX4 $T=1359600 1440880 0 180 $X=1356300 $Y=1435440
X1420 5023 4868 1 3 BUFX4 $T=1550340 1571920 0 0 $X=1550338 $Y=1571518
X1421 5474 5115 1 3 BUFX4 $T=1648020 1521520 0 180 $X=1644720 $Y=1516080
X1422 5909 573 1 3 BUFX4 $T=1942380 1582000 1 0 $X=1942378 $Y=1576560
X1423 602 597 1 3 BUFX4 $T=2033460 1602160 1 180 $X=2030160 $Y=1601758
X1424 4040 315 1 3 317 NAND2BX4 $T=1296900 1481200 0 0 $X=1296898 $Y=1480798
X1425 2577 4416 1 3 4414 NAND2BX4 $T=1387980 1501360 1 0 $X=1387978 $Y=1495920
X1426 2518 4479 1 3 4478 NAND2BX4 $T=1406460 1521520 1 180 $X=1401180 $Y=1521118
X1427 4749 4686 1 3 239 NAND2BX4 $T=1474440 1602160 0 180 $X=1469160 $Y=1596720
X1428 3498 219 161 3 3481 159 1 3476 AOI32X1 $T=1157640 1461040 0 180 $X=1153020 $Y=1455600
X1429 467 6014 6016 3 488 6018 1 6030 AOI32X1 $T=1788600 1511440 1 0 $X=1788598 $Y=1506000
X1430 6125 6097 504 3 6100 498 1 6140 AOI32X1 $T=1815000 1501360 1 0 $X=1814998 $Y=1495920
X1431 6424 6414 553 3 6422 550 1 555 AOI32X1 $T=1895520 1440880 0 0 $X=1895518 $Y=1440478
X1432 9046 9084 742 3 9103 9102 1 744 AOI32X1 $T=2570700 1450960 0 0 $X=2570698 $Y=1450558
X1433 522 6226 1 6228 6233 526 527 3 5946 OAI33X1 $T=1840740 1471120 0 0 $X=1840738 $Y=1470718
X1434 6214 543 1 6394 6398 546 548 3 5945 OAI33X1 $T=1882320 1440880 1 0 $X=1882318 $Y=1435440
X1435 5194 5103 5022 3 1 415 OR3XL $T=1573440 1541680 0 0 $X=1573438 $Y=1541278
X1436 422 5226 5273 3 1 5393 OR3XL $T=1605120 1612240 0 0 $X=1605118 $Y=1611838
X1437 5025 5103 5194 3 1 398 OR3XL $T=1607760 1541680 0 0 $X=1607758 $Y=1541278
X1438 527 526 6285 3 1 6228 OR3XL $T=1851300 1471120 1 180 $X=1848000 $Y=1470718
X1439 548 546 552 3 1 6394 OR3XL $T=1897500 1440880 0 180 $X=1894200 $Y=1435440
X1440 2619 105 1 2619 121 2620 3 OAI22XL $T=944460 1582000 1 0 $X=944458 $Y=1576560
X1441 2690 94 1 2690 2689 2729 3 OAI22XL $T=954360 1561840 0 0 $X=954358 $Y=1561438
X1442 5388 5391 5253 1 396 3 433 OAI31X1 $T=1624260 1491280 1 0 $X=1624258 $Y=1485840
X1443 3 6029 492 6034 493 6038 1 NOR4X1 $T=1793880 1430800 0 0 $X=1793878 $Y=1430398
X1444 2949 1 159 3 161 2973 NAND3XL $T=1018380 1501360 1 0 $X=1018378 $Y=1495920
X1445 436 1 439 3 5246 5508 NAND3XL $T=1658580 1440880 0 180 $X=1655940 $Y=1435440
X1446 5256 403 3 328 5326 1 425 5321 AOI221XL $T=1605780 1582000 1 0 $X=1605778 $Y=1576560
X1447 382 383 381 1 379 3 OAI2BB1XL $T=1508760 1511440 1 180 $X=1505460 $Y=1511038
X1448 254 256 1 258 213 3 250 260 3603 OAI222X1 $T=1209120 1602160 0 0 $X=1209118 $Y=1601758
X1449 322 4139 1 258 227 3 329 260 327 OAI222X1 $T=1332540 1602160 0 180 $X=1326600 $Y=1596720
X1450 5204 5112 1 419 5164 3 5180 5147 5045 OAI222X1 $T=1574100 1511440 0 180 $X=1568160 $Y=1506000
X1451 726 9097 1 9080 739 3 740 9079 9095 OAI222X1 $T=2574660 1582000 1 180 $X=2568720 $Y=1581598
X1452 110 1 105 3 CLKINVX8 $T=881100 1571920 0 0 $X=881098 $Y=1571518
X1453 4721 1 3883 3 CLKINVX8 $T=1461240 1501360 0 0 $X=1461238 $Y=1500958
X1454 392 1 5241 3 CLKINVX8 $T=1579380 1561840 0 0 $X=1579378 $Y=1561438
X1455 5382 1 431 3 CLKINVX8 $T=1625580 1592080 0 0 $X=1625578 $Y=1591678
X1456 5299 1 5534 3 CLKINVX8 $T=1656600 1551760 0 180 $X=1652640 $Y=1546320
X1457 5625 1 4747 3 CLKINVX8 $T=1686960 1491280 1 0 $X=1686958 $Y=1485840
X1458 562 1 561 3 CLKINVX8 $T=1940400 1501360 0 0 $X=1940398 $Y=1500958
X1459 5153 3 5063 1 5113 403 NOR3X1 $T=1566180 1531600 1 0 $X=1566178 $Y=1526160
X1460 424 3 407 1 4744 5134 NOR3X1 $T=1602480 1582000 1 180 $X=1599840 $Y=1581598
X1461 5355 3 407 1 404 5256 NOR3X1 $T=1620960 1582000 0 0 $X=1620958 $Y=1581598
X1462 434 3 407 1 404 5326 NOR3X1 $T=1631520 1561840 1 180 $X=1628880 $Y=1561438
X1463 5498 3 436 1 439 5500 NOR3X1 $T=1653960 1501360 1 0 $X=1653958 $Y=1495920
X1464 4054 4041 3 1 3923 NOR2BX4 $T=1298880 1511440 1 180 $X=1293600 $Y=1511038
X1465 410 5236 3 1 383 NOR2BX4 $T=1580040 1561840 1 0 $X=1580038 $Y=1556400
X1466 5246 5461 3 1 437 NOR2BX4 $T=1653300 1450960 1 180 $X=1648020 $Y=1450558
X1467 6941 6946 3 1 6960 NOR2BX4 $T=2026200 1481200 1 0 $X=2026198 $Y=1475760
X1468 2569 105 121 1 2569 3 121 105 2578 OAI222XL $T=929280 1582000 1 0 $X=929278 $Y=1576560
X1469 2578 2304 39 1 2578 3 2304 39 2683 OAI222XL $T=931920 1561840 0 0 $X=931918 $Y=1561438
X1470 2683 94 94 1 2689 3 2683 2689 2702 OAI222XL $T=951060 1561840 1 0 $X=951058 $Y=1556400
X1471 2702 2728 40 1 2702 3 2728 40 2771 OAI222XL $T=960960 1551760 0 0 $X=960958 $Y=1551358
X1472 2936 99 2936 1 2905 3 2905 99 2950 OAI222XL $T=1013100 1561840 0 0 $X=1013098 $Y=1561438
X1473 90 2950 139 1 2950 3 90 139 2986 OAI222XL $T=1025640 1571920 1 0 $X=1025638 $Y=1566480
X1474 1770 215 211 1 208 3 90 202 3355 OAI222XL $T=1145100 1592080 1 180 $X=1139820 $Y=1591678
X1475 215 2689 213 1 212 3 202 103 3340 OAI222XL $T=1146420 1602160 0 180 $X=1141140 $Y=1596720
X1476 72 215 220 1 212 3 202 3261 3178 OAI222XL $T=1158960 1602160 0 180 $X=1153680 $Y=1596720
X1477 2905 229 227 1 212 3 3493 202 3320 OAI222XL $T=1177440 1602160 0 180 $X=1172160 $Y=1596720
X1478 215 196 243 1 208 3 202 2304 3614 OAI222XL $T=1193280 1602160 0 180 $X=1188000 $Y=1596720
X1479 215 3551 255 1 208 3 202 3604 3679 OAI222XL $T=1203840 1592080 0 0 $X=1203838 $Y=1591678
X1480 251 256 258 1 259 3 248 260 3698 OAI222XL $T=1205160 1612240 0 0 $X=1205158 $Y=1611838
X1481 291 256 258 1 255 3 302 260 3965 OAI222XL $T=1274460 1602160 1 0 $X=1274458 $Y=1596720
X1482 229 2966 316 1 208 3 318 2213 3941 OAI222XL $T=1298220 1592080 0 0 $X=1298218 $Y=1591678
X1483 310 4139 258 1 316 3 307 260 4175 OAI222XL $T=1330560 1592080 0 0 $X=1330558 $Y=1591678
X1484 323 4139 258 1 220 3 321 260 4238 OAI222XL $T=1348380 1612240 0 180 $X=1343100 $Y=1606800
X1485 245 338 258 1 211 3 330 260 4319 OAI222XL $T=1354320 1592080 0 0 $X=1354318 $Y=1591678
X1486 5022 5100 5101 1 5070 3 5110 5112 5107 OAI222XL $T=1550340 1501360 0 0 $X=1550338 $Y=1500958
X1487 5112 5227 5113 1 5132 3 5164 5195 5203 OAI222XL $T=1578060 1501360 0 180 $X=1572780 $Y=1495920
X1488 5115 5253 5164 1 5329 3 5112 5349 5323 OAI222XL $T=1607760 1501360 0 0 $X=1607758 $Y=1500958
X1489 114 2478 1 3 2496 AND2X4 $T=905520 1571920 0 0 $X=905518 $Y=1571518
X1490 5517 5559 1 3 5568 AND2X4 $T=1667820 1592080 1 0 $X=1667818 $Y=1586640
X1491 5693 457 455 1 3 5700 MX2X1 $T=1699500 1582000 0 0 $X=1699498 $Y=1581598
X1492 5693 458 459 1 3 5756 MX2X1 $T=1704780 1612240 1 0 $X=1704778 $Y=1606800
X1493 3980 3 1 206 BUFX8 $T=1279740 1551760 0 180 $X=1273800 $Y=1546320
X1494 388 3 1 4745 BUFX8 $T=1527900 1602160 1 180 $X=1521960 $Y=1601758
X1495 392 3 1 5208 BUFX8 $T=1568820 1602160 0 0 $X=1568818 $Y=1601758
X1496 5241 3 1 4723 BUFX8 $T=1585320 1561840 1 0 $X=1585318 $Y=1556400
X1497 6758 3 1 6781 BUFX8 $T=1981980 1481200 1 0 $X=1981978 $Y=1475760
X1498 2728 40 1 124 3 2729 2726 OAI211XL $T=966240 1571920 0 180 $X=962280 $Y=1566480
X1499 129 128 40 3220 182 3 1 3179 SDFFRHQX1 $T=1095600 1612240 1 180 $X=1079100 $Y=1611838
X1500 129 128 105 3342 122 3 1 3288 SDFFRHQX1 $T=1124640 1612240 0 180 $X=1108140 $Y=1606800
X1501 332 464 553 6538 541 3 1 529 SDFFRHQX1 $T=1916640 1551760 0 0 $X=1916638 $Y=1551358
X1502 332 547 594 6658 541 3 1 6798 SDFFRHQX1 $T=2007060 1582000 1 180 $X=1990560 $Y=1581598
X1503 129 128 47 2760 122 2708 1 3 SDFFRHQX2 $T=975480 1602160 1 180 $X=955680 $Y=1601758
X1504 332 464 478 6331 541 531 1 3 SDFFRHQX2 $T=1861200 1561840 0 0 $X=1861198 $Y=1561438
X1505 3838 41 1 3 BUFX12 $T=1240800 1612240 1 180 $X=1234200 $Y=1611838
X1506 3881 199 1 3 BUFX12 $T=1250700 1511440 0 0 $X=1250698 $Y=1511038
X1507 3923 197 1 3 BUFX12 $T=1257960 1481200 1 0 $X=1257958 $Y=1475760
X1508 3955 207 1 3 BUFX12 $T=1271820 1511440 1 180 $X=1265220 $Y=1511038
X1509 5241 5255 1 3 BUFX12 $T=1584660 1551760 0 0 $X=1584658 $Y=1551358
X1510 5896 471 1 3 BUFX12 $T=1752960 1612240 1 0 $X=1752958 $Y=1606800
X1511 129 139 128 3178 122 3 1 130 SDFFRHQX4 $T=1075140 1571920 0 0 $X=1075138 $Y=1571518
X1512 129 218 241 3614 232 3 1 104 SDFFRHQX4 $T=1198560 1561840 0 180 $X=1174140 $Y=1556400
X1513 129 272 128 3941 182 3 1 108 SDFFRHQX4 $T=1269840 1571920 1 180 $X=1245420 $Y=1571518
X1514 1770 42 52 3 1781 1782 1 AOI2BB2XL $T=716100 1511440 0 0 $X=716098 $Y=1511038
X1515 1770 224 225 3 226 3557 1 AOI2BB2XL $T=1171500 1592080 0 0 $X=1171498 $Y=1591678
X1516 121 239 240 3 237 3613 1 AOI2BB2XL $T=1187340 1612240 0 0 $X=1187338 $Y=1611838
X1517 3551 224 270 3 268 3777 1 AOI2BB2XL $T=1222320 1592080 0 0 $X=1222318 $Y=1591678
X1518 2905 239 289 3 237 3876 1 AOI2BB2XL $T=1244760 1602160 0 0 $X=1244758 $Y=1601758
X1519 2966 239 306 3 268 4012 1 AOI2BB2XL $T=1291620 1602160 0 180 $X=1287000 $Y=1596720
X1520 477 398 427 3 478 5990 1 AOI2BB2XL $T=1778040 1592080 1 0 $X=1778038 $Y=1586640
X1521 503 415 414 3 501 6116 1 AOI2BB2XL $T=1814340 1582000 1 180 $X=1809720 $Y=1581598
X1522 520 415 414 3 6157 6158 1 AOI2BB2XL $T=1824900 1582000 1 180 $X=1820280 $Y=1581598
X1523 242 254 250 247 3624 2760 3 1 OAI221X4 $T=1203840 1612240 0 180 $X=1196580 $Y=1606800
X1524 242 310 307 304 4012 2749 3 1 OAI221X4 $T=1291620 1592080 1 180 $X=1284360 $Y=1591678
X1525 129 128 49 3230 122 1770 139 1 3 SDFFRX4 $T=1098240 1582000 1 180 $X=1075140 $Y=1581598
X1526 129 241 214 3679 232 3604 80 1 3 SDFFRX4 $T=1199220 1561840 0 0 $X=1199218 $Y=1561438
X1527 129 241 192 280 232 284 101 1 3 SDFFRX4 $T=1234200 1511440 1 0 $X=1234198 $Y=1506000
X1528 409 1 416 5324 5355 5315 3 NAND4X1 $T=1613700 1592080 1 0 $X=1613698 $Y=1586640
X1529 407 1 5198 414 5208 5559 3 NAND4X1 $T=1640100 1582000 0 0 $X=1640098 $Y=1581598
X1530 198 1 3 3413 BUFXL $T=1144440 1582000 0 0 $X=1144438 $Y=1581598
X1531 198 1 3 3514 BUFXL $T=1164240 1551760 0 0 $X=1164238 $Y=1551358
X1532 392 1 3 5064 BUFXL $T=1549680 1592080 1 0 $X=1549678 $Y=1586640
X1533 5400 1 3 5407 BUFXL $T=1627560 1612240 1 0 $X=1627558 $Y=1606800
X1534 5208 1 3 5513 BUFXL $T=1644720 1582000 0 0 $X=1644718 $Y=1581598
X1535 4152 4166 4131 3 4204 4155 1 AOI31X2 $T=1325280 1531600 1 0 $X=1325278 $Y=1526160
X1536 4233 4212 4224 3 4204 4205 1 AOI31X2 $T=1343760 1531600 0 180 $X=1337820 $Y=1526160
X1537 4249 4248 4120 3 4204 4293 1 AOI31X2 $T=1349700 1541680 1 0 $X=1349698 $Y=1536240
X1538 4304 4302 4288 3 4204 4292 1 AOI31X2 $T=1358280 1521520 1 180 $X=1352340 $Y=1521118
X1539 6158 505 508 3 487 507 1 AOI31X2 $T=1818300 1592080 0 180 $X=1812360 $Y=1586640
X1540 5293 1 421 410 3 5319 NAND3X4 $T=1599180 1521520 0 0 $X=1599178 $Y=1521118
X1541 6345 1 6209 6356 3 6331 NAND3BX1 $T=1869120 1592080 0 0 $X=1869118 $Y=1591678
X1542 470 1 5894 3 CLKINVX2 $T=1756260 1551760 1 180 $X=1754280 $Y=1551358
X1543 5401 5404 5406 5400 3 1 5382 NAND4X4 $T=1620960 1602160 1 0 $X=1620958 $Y=1596720
X1544 6498 542 545 561 3 1 6509 NAND4X4 $T=1914000 1501360 0 180 $X=1902780 $Y=1495920
X1545 414 5129 3 5268 1 5201 5272 AOI211XL $T=1591260 1561840 1 0 $X=1591258 $Y=1556400
X1546 510 503 1 500 289 6124 3 AOI2BB2X2 $T=1815660 1602160 0 180 $X=1809720 $Y=1596720
X1547 189 186 190 3 1 3190 ADDHX1 $T=1105500 1450960 1 180 $X=1097580 $Y=1450558
X1548 426 1 3 428 CLKBUFX20 $T=1605780 1440880 0 0 $X=1605778 $Y=1440478
X1549 5208 5207 397 5226 377 3 1 OAI31X4 $T=1577400 1612240 0 0 $X=1577398 $Y=1611838
X1550 4155 4530 352 3 4543 4529 1 NAND4BBX1 $T=1417020 1471120 1 0 $X=1417018 $Y=1465680
X1551 4831 4835 1 4841 374 3 NAND3BX4 $T=1491600 1592080 0 0 $X=1491598 $Y=1591678
X1552 5113 3 5063 1 5103 5001 NOR3XL $T=1552980 1531600 0 180 $X=1550340 $Y=1526160
X1553 5103 3 5150 1 5022 391 NOR3XL $T=1558260 1541680 1 180 $X=1555620 $Y=1541278
X1554 5494 3 436 1 5236 5510 NOR3XL $T=1651980 1471120 1 180 $X=1649340 $Y=1470718
X1555 332 241 5063 5203 234 5113 1 3 5200 SDFFSXL $T=1574100 1461040 1 0 $X=1574098 $Y=1455600
X1556 410 5246 1 3 CLKBUFX4 $T=1582680 1541680 0 0 $X=1582678 $Y=1541278
X1557 5272 1 5330 5038 5149 5260 3 NAND4XL $T=1594560 1551760 1 180 $X=1591260 $Y=1551358
X1558 5534 1 5536 5537 5474 5543 3 NAND4XL $T=1661220 1551760 1 0 $X=1661218 $Y=1546320
X1559 5579 1 441 5508 5533 5543 3 NAND4XL $T=1667160 1440880 0 180 $X=1663860 $Y=1435440
X1560 5329 5197 3 5327 5129 414 5361 5349 1 AOI222XL $T=1613040 1511440 0 0 $X=1613038 $Y=1511038
X1561 5404 1 3 5420 BUFX1 $T=1632180 1592080 0 0 $X=1632178 $Y=1591678
X1562 389 5051 5023 1 5239 5404 3 AOI2BB2X4 $T=1632180 1602160 1 0 $X=1632178 $Y=1596720
X1563 388 398 5208 1 5207 5406 3 AOI2BB2X4 $T=1650000 1592080 0 0 $X=1649998 $Y=1591678
X1564 388 398 5208 1 5207 5517 3 AOI2BB2X4 $T=1650000 1602160 1 0 $X=1649998 $Y=1596720
X1565 562 528 6541 559 563 1 3 OR4X4 $T=1921260 1501360 0 0 $X=1921258 $Y=1500958
X1566 7856 7859 7810 7825 1 3 7075 OAI2BB2XL $T=2251260 1541680 1 180 $X=2246640 $Y=1541278
.ENDS
***************************************
.SUBCKT ADDHX2 B S A VDD VSS CO
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRX1 CK SE SI D RN QN VDD VSS Q
** N=11 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4BX4 AN B C D VDD VSS Y
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_58 2 4 42 43 44 45 46 47 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 86 87 88 89 92 93 95 96 98 99 100 103 104 105 106 107
+ 108 109 111 112 113 115 116 117 118 119 123 124 125 126 127 128 129 130 131 132
+ 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152
+ 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 174
+ 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 191 192 193 194 195
+ 196 197 198 199 200 202 203 205 206 207 208 209 210 211 213 214 215 216 217 218
+ 219 221 222 223 224 225 226 227 228 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 355 356 357 358 359 360 361
+ 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381
+ 382 383 384 385 386 387 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 413 414 416 417 418 420 421 422 423 424 426
+ 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446
+ 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466
+ 467 468 469 470 471 472 473 475 476 477 478 479 480 481 482 484 485 487 488 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 524 525 527 528 529 530 531 532
+ 534 535 536 537 538 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554
+ 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574
+ 576 577 578 580 581 583 584 585 587 588 589 590 592 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 625 626 627 628 630 631 632 633 634 636 637 639 641 643 644 646 647
+ 649 650 651 652 653 654 655 656 657 658 659 660 661 662 663 664 665 667 668 669
+ 671 672 674 675 676 677 678 679 680 681 682 683 684 685 686 687 688 689 690 691
+ 692 693 694 695 697 698 699 700 701 702 704 705 707 708 709 710 711 712 713 714
+ 715 716 717 719 720 722 724 725 726 728 730 732 733 734 735 736 737 778 779 780
+ 781 782 783 784 785 786 787 788 789 1652 1653
** N=35507 EP=651 IP=13281 FDC=0
X0 53 2 54 4 1886 NAND2X1 $T=716100 2065840 0 0 $X=716098 $Y=2065438
X1 59 2 54 4 1924 NAND2X1 $T=726000 2075920 0 180 $X=724020 $Y=2070480
X2 2057 2 2060 4 69 NAND2X1 $T=751740 2217040 1 0 $X=751738 $Y=2211600
X3 2097 2 2093 4 74 NAND2X1 $T=762960 2196880 1 180 $X=760980 $Y=2196478
X4 2134 2 2136 4 80 NAND2X1 $T=776160 2186800 1 180 $X=774180 $Y=2186398
X5 2299 2 2319 4 2337 NAND2X1 $T=813120 2206960 1 0 $X=813118 $Y=2201520
X6 2382 2 2296 4 2359 NAND2X1 $T=817740 2186800 1 180 $X=815760 $Y=2186398
X7 2565 2 2560 4 2588 NAND2X1 $T=862620 2146480 1 0 $X=862618 $Y=2141040
X8 2636 2 2614 4 2633 NAND2X1 $T=875160 2136400 0 180 $X=873180 $Y=2130960
X9 2603 2 2630 4 2667 NAND2X1 $T=878460 2146480 1 0 $X=878458 $Y=2141040
X10 2610 2 2590 4 2636 NAND2X1 $T=883740 2116240 1 0 $X=883738 $Y=2110800
X11 2707 2 2665 4 2708 NAND2X1 $T=893640 2116240 0 180 $X=891660 $Y=2110800
X12 2716 2 2614 4 2721 NAND2X1 $T=893640 2136400 1 0 $X=893638 $Y=2130960
X13 2801 2 2789 4 2839 NAND2X1 $T=914760 2075920 0 0 $X=914758 $Y=2075518
X14 2843 2 2841 4 2844 NAND2X1 $T=917400 2086000 1 180 $X=915420 $Y=2085598
X15 2913 2 2710 4 2863 NAND2X1 $T=925980 2206960 1 180 $X=924000 $Y=2206558
X16 2843 2 2834 4 2906 NAND2X1 $T=926640 2086000 1 0 $X=926638 $Y=2080560
X17 2711 2 2830 4 2928 NAND2X1 $T=927960 2055760 0 0 $X=927958 $Y=2055358
X18 2928 2 2843 4 2945 NAND2X1 $T=935220 2086000 1 180 $X=933240 $Y=2085598
X19 2989 2 2959 4 2956 NAND2X1 $T=939840 2166640 0 180 $X=937860 $Y=2161200
X20 95 2 71 4 3066 NAND2X1 $T=941160 2025520 0 0 $X=941158 $Y=2025118
X21 2421 2 55 4 3059 NAND2X1 $T=943800 2045680 0 0 $X=943798 $Y=2045278
X22 3066 2 3064 4 3106 NAND2X1 $T=957000 2025520 1 0 $X=956998 $Y=2020080
X23 3058 2 3085 4 3114 NAND2X1 $T=957000 2196880 1 0 $X=956998 $Y=2191440
X24 93 2 51 4 3110 NAND2X1 $T=964260 2055760 1 180 $X=962280 $Y=2055358
X25 3146 2 3120 4 3118 NAND2X1 $T=964920 2136400 1 180 $X=962940 $Y=2135998
X26 3136 2 3119 4 3120 NAND2X1 $T=965580 2126320 1 180 $X=963600 $Y=2125918
X27 3117 2 3184 4 116 NAND2X1 $T=969540 2186800 0 0 $X=969538 $Y=2186398
X28 3207 2 2938 4 3159 NAND2X1 $T=972180 2025520 0 180 $X=970200 $Y=2020080
X29 3187 2 3138 4 3146 NAND2X1 $T=972180 2126320 0 180 $X=970200 $Y=2120880
X30 3199 2 3186 4 3200 NAND2X1 $T=978780 2065840 1 180 $X=976800 $Y=2065438
X31 3230 2 2977 4 3195 NAND2X1 $T=983400 2106160 0 180 $X=981420 $Y=2100720
X32 3333 2 3329 4 3327 NAND2X1 $T=1001880 2025520 1 180 $X=999900 $Y=2025118
X33 3444 2 3412 4 3432 NAND2X1 $T=1017720 2156560 0 180 $X=1015740 $Y=2151120
X34 3416 2 3122 4 3411 NAND2X1 $T=1019040 2035600 0 180 $X=1017060 $Y=2030160
X35 3411 2 3435 4 3464 NAND2X1 $T=1022340 2065840 1 0 $X=1022338 $Y=2060400
X36 3481 2 3255 4 3438 NAND2X1 $T=1024980 2055760 0 180 $X=1023000 $Y=2050320
X37 3471 2 3431 4 3479 NAND2X1 $T=1030260 2116240 0 0 $X=1030258 $Y=2115838
X38 3418 2 3482 4 3364 NAND2X1 $T=1030260 2166640 0 0 $X=1030258 $Y=2166238
X39 125 2 124 4 3508 NAND2X1 $T=1037520 1995280 0 180 $X=1035540 $Y=1989840
X40 3553 2 3562 4 3359 NAND2X1 $T=1046760 2196880 1 0 $X=1046758 $Y=2191440
X41 3569 2 3564 4 3494 NAND2X1 $T=1048740 2096080 0 180 $X=1046760 $Y=2090640
X42 3659 2 3658 4 3660 NAND2X1 $T=1063260 2075920 1 180 $X=1061280 $Y=2075518
X43 131 2 128 4 3461 NAND2X1 $T=1065240 2005360 1 0 $X=1065238 $Y=1999920
X44 137 2 3639 4 3640 NAND2X1 $T=1068540 2035600 0 180 $X=1066560 $Y=2030160
X45 3698 2 3626 4 3566 NAND2X1 $T=1071840 2106160 1 0 $X=1071838 $Y=2100720
X46 3464 2 3703 4 3705 NAND2X1 $T=1073160 2065840 0 0 $X=1073158 $Y=2065438
X47 3769 2 3256 4 3781 NAND2X1 $T=1090320 2065840 1 0 $X=1090318 $Y=2060400
X48 3783 2 148 4 3724 NAND2X1 $T=1092300 2025520 0 180 $X=1090320 $Y=2020080
X49 3815 2 152 4 3861 NAND2X1 $T=1106160 2025520 1 0 $X=1106158 $Y=2020080
X50 3956 2 95 4 3915 NAND2X1 $T=1122000 2055760 0 180 $X=1120020 $Y=2050320
X51 3794 2 163 4 168 NAND2X1 $T=1121340 1995280 0 0 $X=1121338 $Y=1994878
X52 140 2 3958 4 3917 NAND2X1 $T=1131900 2015440 0 0 $X=1131898 $Y=2015038
X53 4321 2 203 4 4443 NAND2X1 $T=1228920 2015440 0 0 $X=1228918 $Y=2015038
X54 4486 2 4480 4 226 NAND2X1 $T=1238160 2227120 0 180 $X=1236180 $Y=2221680
X55 4599 2 195 4 4507 NAND2X1 $T=1246740 2075920 1 180 $X=1244760 $Y=2075518
X56 4535 2 4505 4 4659 NAND2X1 $T=1256640 2096080 0 0 $X=1256638 $Y=2095678
X57 244 2 252 4 4735 NAND2X1 $T=1288980 2106160 0 0 $X=1288978 $Y=2105758
X58 4765 2 4786 4 4741 NAND2X1 $T=1296900 2045680 0 0 $X=1296898 $Y=2045278
X59 264 2 3140 4 4891 NAND2X1 $T=1312080 2217040 0 180 $X=1310100 $Y=2211600
X60 4891 2 4908 4 5108 NAND2X1 $T=1323300 2206960 0 0 $X=1323298 $Y=2206558
X61 4949 2 4932 4 4890 NAND2X1 $T=1325280 2075920 1 180 $X=1323300 $Y=2075518
X62 3188 2 271 4 4995 NAND2X1 $T=1333200 2196880 0 180 $X=1331220 $Y=2191440
X63 4851 2 4968 4 4949 NAND2X1 $T=1331880 2096080 0 0 $X=1331878 $Y=2095678
X64 4994 2 4908 4 5004 NAND2X1 $T=1339140 2206960 1 180 $X=1337160 $Y=2206558
X65 4995 2 4994 4 5026 NAND2X1 $T=1338480 2196880 1 0 $X=1338478 $Y=2191440
X66 4998 2 4954 4 5012 NAND2X1 $T=1340460 2065840 1 180 $X=1338480 $Y=2065438
X67 5002 2 4998 4 4972 NAND2X1 $T=1341780 2055760 1 180 $X=1339800 $Y=2055358
X68 3337 2 275 4 5019 NAND2X1 $T=1343100 2156560 1 180 $X=1341120 $Y=2156158
X69 5076 2 5040 4 5002 NAND2X1 $T=1349700 2055760 1 180 $X=1347720 $Y=2055358
X70 5003 2 5074 4 4978 NAND2X1 $T=1350360 2086000 0 0 $X=1350358 $Y=2085598
X71 4980 2 4996 4 5038 NAND2X1 $T=1356960 2005360 1 0 $X=1356958 $Y=1999920
X72 5096 2 5123 4 5126 NAND2X1 $T=1362240 2005360 0 0 $X=1362238 $Y=2004958
X73 3392 2 286 4 5192 NAND2X1 $T=1375440 2096080 1 0 $X=1375438 $Y=2090640
X74 5192 2 5234 4 5248 NAND2X1 $T=1387980 2106160 1 0 $X=1387978 $Y=2100720
X75 3387 2 5323 4 5343 NAND2X1 $T=1402500 2075920 1 0 $X=1402498 $Y=2070480
X76 5343 2 5366 4 5437 NAND2X1 $T=1424940 2075920 1 0 $X=1424938 $Y=2070480
X77 3702 2 345 4 5886 NAND2X1 $T=1516680 2086000 1 0 $X=1516678 $Y=2080560
X78 5889 2 3667 4 5982 NAND2X1 $T=1537140 2096080 0 0 $X=1537138 $Y=2095678
X79 5982 2 5961 4 6051 NAND2X1 $T=1550340 2086000 0 0 $X=1550338 $Y=2085598
X80 6058 2 4108 4 6059 NAND2X1 $T=1564860 2075920 1 0 $X=1564858 $Y=2070480
X81 6191 2 4086 4 6257 NAND2X1 $T=1604460 2045680 0 0 $X=1604458 $Y=2045278
X82 6270 2 4637 4 6249 NAND2X1 $T=1609740 2015440 1 0 $X=1609738 $Y=2010000
X83 6338 2 4742 4 6335 NAND2X1 $T=1625580 2005360 1 180 $X=1623600 $Y=2004958
X84 6345 2 6440 4 6425 NAND2X1 $T=1645380 2005360 0 0 $X=1645378 $Y=2004958
X85 6338 2 6440 4 6517 NAND2X1 $T=1664520 2005360 0 0 $X=1664518 $Y=2004958
X86 6591 2 6440 4 416 NAND2X1 $T=1693560 1995280 1 0 $X=1693558 $Y=1989840
X87 6723 2 6057 4 6715 NAND2X1 $T=1704120 2075920 0 180 $X=1702140 $Y=2070480
X88 6720 2 417 4 6697 NAND2X1 $T=1706760 2005360 0 180 $X=1704780 $Y=1999920
X89 400 2 409 4 6714 NAND2X1 $T=1706100 2055760 0 0 $X=1706098 $Y=2055358
X90 6807 2 6080 4 6759 NAND2X1 $T=1731840 2015440 0 0 $X=1731838 $Y=2015038
X91 6768 2 432 4 6850 NAND2X1 $T=1736460 2065840 1 0 $X=1736458 $Y=2060400
X92 438 2 409 4 442 NAND2X1 $T=1746360 2035600 0 180 $X=1744380 $Y=2030160
X93 6944 2 5741 4 6869 NAND2X1 $T=1749000 2075920 0 180 $X=1747020 $Y=2070480
X94 6986 2 6964 4 6990 NAND2X1 $T=1764180 2096080 0 180 $X=1762200 $Y=2090640
X95 7030 2 5362 4 6986 NAND2X1 $T=1770120 2106160 0 180 $X=1768140 $Y=2100720
X96 7026 2 457 4 6989 NAND2X1 $T=1780680 2035600 0 0 $X=1780678 $Y=2035198
X97 7080 2 465 4 7047 NAND2X1 $T=1793220 2065840 0 180 $X=1791240 $Y=2060400
X98 7168 2 469 4 7101 NAND2X1 $T=1802460 2045680 1 180 $X=1800480 $Y=2045278
X99 7194 2 7170 4 7169 NAND2X1 $T=1804440 2106160 1 180 $X=1802460 $Y=2105758
X100 7188 2 5260 4 7166 NAND2X1 $T=1807740 2126320 0 180 $X=1805760 $Y=2120880
X101 7189 2 470 4 7059 NAND2X1 $T=1808400 2015440 0 0 $X=1808398 $Y=2015038
X102 7255 2 479 4 7208 NAND2X1 $T=1822260 2005360 0 180 $X=1820280 $Y=1999920
X103 7256 2 7252 4 478 NAND2X1 $T=1822260 2025520 1 180 $X=1820280 $Y=2025118
X104 7261 2 5149 4 7257 NAND2X1 $T=1822260 2075920 1 180 $X=1820280 $Y=2075518
X105 7297 2 7260 4 7256 NAND2X1 $T=1824240 2035600 1 180 $X=1822260 $Y=2035198
X106 7300 2 7296 4 7252 NAND2X1 $T=1832160 2025520 1 180 $X=1830180 $Y=2025118
X107 7433 2 487 4 7354 NAND2X1 $T=1843380 2075920 1 180 $X=1841400 $Y=2075518
X108 7471 2 5152 4 7378 NAND2X1 $T=1857240 2106160 1 180 $X=1855260 $Y=2105758
X109 7455 2 490 4 7374 NAND2X1 $T=1857240 2025520 1 0 $X=1857238 $Y=2020080
X110 7587 2 495 4 7603 NAND2X1 $T=1888260 2065840 0 0 $X=1888258 $Y=2065438
X111 502 2 497 4 7592 NAND2X1 $T=1891560 2126320 1 180 $X=1889580 $Y=2125918
X112 509 2 7745 4 7790 NAND2X1 $T=1917300 2196880 0 0 $X=1917298 $Y=2196478
X113 514 2 516 4 7788 NAND2X1 $T=1935120 2055760 0 0 $X=1935118 $Y=2055358
X114 7939 2 528 4 7907 NAND2X1 $T=1959540 2126320 0 0 $X=1959538 $Y=2125918
X115 8024 2 541 4 8057 NAND2X1 $T=1978020 2116240 0 0 $X=1978018 $Y=2115838
X116 8188 2 8210 4 8235 NAND2X1 $T=2009700 2176720 1 0 $X=2009698 $Y=2171280
X117 8258 2 8236 4 8194 NAND2X1 $T=2013000 2015440 1 180 $X=2011020 $Y=2015038
X118 8263 2 564 4 8188 NAND2X1 $T=2020260 2176720 1 180 $X=2018280 $Y=2176318
X119 561 2 563 4 8258 NAND2X1 $T=2019600 2005360 1 0 $X=2019598 $Y=1999920
X120 8305 2 8282 4 8288 NAND2X1 $T=2023560 2126320 0 180 $X=2021580 $Y=2120880
X121 565 2 8291 4 8305 NAND2X1 $T=2028840 2106160 0 180 $X=2026860 $Y=2100720
X122 573 2 8323 4 8281 NAND2X1 $T=2032800 2025520 0 180 $X=2030820 $Y=2020080
X123 8329 2 570 4 8312 NAND2X1 $T=2033460 2196880 0 0 $X=2033458 $Y=2196478
X124 8405 2 578 4 8439 NAND2X1 $T=2055240 2206960 0 0 $X=2055238 $Y=2206558
X125 581 2 8454 4 8437 NAND2X1 $T=2058540 2015440 0 180 $X=2056560 $Y=2010000
X126 8438 2 8436 4 8457 NAND2X1 $T=2061180 2136400 0 180 $X=2059200 $Y=2130960
X127 8479 2 8513 4 8493 NAND2X1 $T=2072400 2106160 0 0 $X=2072398 $Y=2105758
X128 8521 2 8512 4 8495 NAND2X1 $T=2074380 2025520 1 180 $X=2072400 $Y=2025118
X129 8516 2 588 4 8555 NAND2X1 $T=2077680 2217040 0 0 $X=2077678 $Y=2216638
X130 590 2 589 4 8510 NAND2X1 $T=2079660 1995280 1 180 $X=2077680 $Y=1994878
X131 8566 2 8591 4 8584 NAND2X1 $T=2089560 2116240 0 0 $X=2089558 $Y=2115838
X132 8672 2 8692 4 8691 NAND2X1 $T=2112660 2126320 0 0 $X=2112658 $Y=2125918
X133 598 2 602 4 8740 NAND2X1 $T=2113980 2005360 1 0 $X=2113978 $Y=1999920
X134 8719 2 8763 4 8724 NAND2X1 $T=2120580 2126320 1 0 $X=2120578 $Y=2120880
X135 8808 2 8829 4 8823 NAND2X1 $T=2136420 2136400 1 0 $X=2136418 $Y=2130960
X136 8812 2 8883 4 8882 NAND2X1 $T=2146980 2146480 1 0 $X=2146978 $Y=2141040
X137 8892 2 8929 4 8890 NAND2X1 $T=2154900 2126320 1 0 $X=2154898 $Y=2120880
X138 619 2 8946 4 8876 NAND2X1 $T=2162820 2015440 0 0 $X=2162818 $Y=2015038
X139 8989 2 620 4 8975 NAND2X1 $T=2169420 2217040 0 0 $X=2169418 $Y=2216638
X140 9015 2 9017 4 9020 NAND2X1 $T=2173380 2146480 1 0 $X=2173378 $Y=2141040
X141 9064 2 623 4 9037 NAND2X1 $T=2179980 2186800 0 180 $X=2178000 $Y=2181360
X142 8990 2 9035 4 9018 NAND2X1 $T=2181300 2116240 0 0 $X=2181298 $Y=2115838
X143 8972 2 9066 4 9023 NAND2X1 $T=2185920 2015440 0 0 $X=2185918 $Y=2015038
X144 9168 2 627 4 9169 NAND2X1 $T=2203740 2217040 1 180 $X=2201760 $Y=2216638
X145 9166 2 9105 4 9098 NAND2X1 $T=2207040 2136400 0 0 $X=2207038 $Y=2135998
X146 9273 2 637 4 9269 NAND2X1 $T=2228820 2005360 1 180 $X=2226840 $Y=2004958
X147 9184 2 9253 4 9281 NAND2X1 $T=2236080 2126320 0 0 $X=2236078 $Y=2125918
X148 9281 2 9320 4 9319 NAND2X1 $T=2238060 2146480 0 0 $X=2238058 $Y=2146078
X149 9322 2 641 4 9342 NAND2X1 $T=2240040 2206960 1 0 $X=2240038 $Y=2201520
X150 9282 2 9356 4 9357 NAND2X1 $T=2245980 2015440 0 0 $X=2245978 $Y=2015038
X151 9344 2 9422 4 9424 NAND2X1 $T=2253900 2217040 1 0 $X=2253898 $Y=2211600
X152 644 2 9245 4 9425 NAND2X1 $T=2255880 2005360 0 180 $X=2253900 $Y=1999920
X153 9488 2 9422 4 9510 NAND2X1 $T=2271060 2217040 1 0 $X=2271058 $Y=2211600
X154 9489 2 650 4 9488 NAND2X1 $T=2273700 2217040 0 0 $X=2273698 $Y=2216638
X155 653 2 651 4 9546 NAND2X1 $T=2288880 1995280 0 180 $X=2286900 $Y=1989840
X156 651 2 654 4 9725 NAND2X1 $T=2306700 1995280 1 0 $X=2306698 $Y=1989840
X157 9514 2 9600 4 9700 NAND2X1 $T=2309340 2126320 0 0 $X=2309338 $Y=2125918
X158 9796 2 9830 4 9735 NAND2X1 $T=2338380 2217040 1 0 $X=2338378 $Y=2211600
X159 9661 2 9809 4 9879 NAND2X1 $T=2343000 2126320 0 0 $X=2342998 $Y=2125918
X160 9859 2 664 4 9796 NAND2X1 $T=2344980 2227120 1 0 $X=2344978 $Y=2221680
X161 9873 2 9861 4 9938 NAND2X1 $T=2347620 2106160 1 180 $X=2345640 $Y=2105758
X162 9918 2 667 4 9930 NAND2X1 $T=2355540 2206960 0 0 $X=2355538 $Y=2206558
X163 9917 2 672 4 9996 NAND2X1 $T=2369400 2217040 1 0 $X=2369398 $Y=2211600
X164 676 2 677 4 10018 NAND2X1 $T=2378640 2227120 0 0 $X=2378638 $Y=2226718
X165 9935 2 10033 4 10136 NAND2X1 $T=2381280 2126320 1 0 $X=2381278 $Y=2120880
X166 10142 2 10074 4 10230 NAND2X1 $T=2417580 2136400 0 0 $X=2417578 $Y=2135998
X167 10201 2 10054 4 10322 NAND2X1 $T=2440020 2116240 0 0 $X=2440018 $Y=2115838
X168 10290 2 10225 4 10325 NAND2X1 $T=2442660 2116240 1 0 $X=2442658 $Y=2110800
X169 10433 2 10432 4 10315 NAND2X1 $T=2461140 2176720 1 180 $X=2459160 $Y=2176318
X170 10462 2 10444 4 10433 NAND2X1 $T=2466420 2186800 1 0 $X=2466418 $Y=2181360
X171 10472 2 10523 4 10522 NAND2X1 $T=2484240 2035600 1 0 $X=2484238 $Y=2030160
X172 10418 2 10518 4 10570 NAND2X1 $T=2489520 2096080 1 0 $X=2489518 $Y=2090640
X173 10560 2 10590 4 10610 NAND2X1 $T=2494800 2136400 1 0 $X=2494798 $Y=2130960
X174 10609 2 10443 4 10683 NAND2X1 $T=2500080 2116240 0 0 $X=2500078 $Y=2115838
X175 10662 2 10685 4 10726 NAND2X1 $T=2514600 2015440 0 0 $X=2514598 $Y=2015038
X176 10682 2 10724 4 704 NAND2X1 $T=2515260 2035600 1 0 $X=2515258 $Y=2030160
X177 10852 2 10787 4 10980 NAND2X1 $T=2536380 2065840 0 0 $X=2536378 $Y=2065438
X178 10937 2 10554 4 10941 NAND2X1 $T=2552220 2086000 0 0 $X=2552218 $Y=2085598
X179 10974 2 10782 4 10982 NAND2X1 $T=2552220 2116240 0 0 $X=2552218 $Y=2115838
X180 10976 2 10977 4 10972 NAND2X1 $T=2553540 2075920 0 0 $X=2553538 $Y=2075518
X181 10989 2 719 4 720 NAND2X1 $T=2556840 2005360 0 180 $X=2554860 $Y=1999920
X182 10977 2 10943 4 11065 NAND2X1 $T=2564760 2096080 0 180 $X=2562780 $Y=2090640
X183 11091 2 10782 4 11043 NAND2X1 $T=2578620 2116240 1 0 $X=2578618 $Y=2110800
X184 11064 2 726 4 728 NAND2X1 $T=2580600 2015440 0 0 $X=2580598 $Y=2015038
X185 11020 2 10844 4 11004 NAND2X1 $T=2589180 2055760 0 0 $X=2589178 $Y=2055358
X186 11155 2 10782 4 11133 NAND2X1 $T=2591160 2116240 0 180 $X=2589180 $Y=2110800
X187 11227 2 733 4 11250 NAND2X1 $T=2604360 2035600 1 0 $X=2604358 $Y=2030160
X188 11250 2 11290 4 737 NAND2X1 $T=2617560 2005360 1 0 $X=2617558 $Y=1999920
X189 2710 4 2 2913 2892 NOR2X4 $T=930600 2206960 0 0 $X=930598 $Y=2206558
X190 3381 4 2 270 4951 NOR2X4 $T=1327920 2146480 1 0 $X=1327918 $Y=2141040
X191 7455 4 2 490 7454 NOR2X4 $T=1861200 2015440 0 180 $X=1856580 $Y=2010000
X192 7471 4 2 5152 7333 NOR2X4 $T=1857240 2116240 0 0 $X=1857238 $Y=2115838
X193 7939 4 2 528 7895 NOR2X4 $T=1955580 2126320 1 180 $X=1950960 $Y=2125918
X194 536 4 2 535 8007 NOR2X4 $T=1966140 2055760 1 0 $X=1966138 $Y=2050320
X195 548 4 2 543 7999 NOR2X4 $T=1987260 2035600 1 0 $X=1987258 $Y=2030160
X196 604 4 2 8742 778 NOR2X4 $T=2115300 2227120 0 0 $X=2115298 $Y=2226718
X197 2397 2 2359 2519 4 NAND2BX1 $T=844140 2227120 1 0 $X=844138 $Y=2221680
X198 2892 2 2863 109 4 NAND2BX1 $T=927960 2227120 1 0 $X=927958 $Y=2221680
X199 3057 2 2956 2986 4 NAND2BX1 $T=948420 2176720 1 180 $X=945780 $Y=2176318
X200 3107 2 3059 3142 4 NAND2BX1 $T=960300 2045680 0 0 $X=960298 $Y=2045278
X201 3145 2 3146 3224 4 NAND2BX1 $T=970200 2136400 0 0 $X=970198 $Y=2135998
X202 3166 2 3195 3206 4 NAND2BX1 $T=981420 2146480 0 0 $X=981418 $Y=2146078
X203 3226 2 3159 3250 4 NAND2BX1 $T=993300 2025520 1 0 $X=993298 $Y=2020080
X204 3231 2 3327 3330 4 NAND2BX1 $T=1001220 2055760 1 0 $X=1001218 $Y=2050320
X205 3362 2 3359 3274 4 NAND2BX1 $T=1006500 2196880 1 180 $X=1003860 $Y=2196478
X206 3389 2 3438 3487 4 NAND2BX1 $T=1026960 2065840 1 0 $X=1026958 $Y=2060400
X207 3541 2 3508 3509 4 NAND2BX1 $T=1037520 2015440 0 180 $X=1034880 $Y=2010000
X208 3560 2 3566 3618 4 NAND2BX1 $T=1056000 2116240 0 180 $X=1053360 $Y=2110800
X209 139 2 132 3787 4 NAND2BX1 $T=1081740 2045680 0 0 $X=1081738 $Y=2045278
X210 3935 2 3917 3962 4 NAND2BX1 $T=1134540 2035600 1 0 $X=1134538 $Y=2030160
X211 3936 2 3915 4027 4 NAND2BX1 $T=1139820 2055760 1 0 $X=1139818 $Y=2050320
X212 252 2 263 4728 4 NAND2BX1 $T=1310760 2106160 1 180 $X=1308120 $Y=2105758
X213 4973 2 4978 4866 4 NAND2BX1 $T=1343760 2086000 1 180 $X=1341120 $Y=2085598
X214 5077 2 5019 5127 4 NAND2BX1 $T=1360920 2136400 0 0 $X=1360918 $Y=2135998
X215 5493 2 328 5397 4 NAND2BX1 $T=1481040 2156560 0 180 $X=1478400 $Y=2151120
X216 5874 2 5886 5966 4 NAND2BX1 $T=1539780 2075920 1 0 $X=1539778 $Y=2070480
X217 6054 2 6059 6117 4 NAND2BX1 $T=1564860 2055760 1 0 $X=1564858 $Y=2050320
X218 6246 2 6249 6299 4 NAND2BX1 $T=1602480 1995280 0 0 $X=1602478 $Y=1994878
X219 6787 2 6759 6758 4 NAND2BX1 $T=1717980 2015440 1 180 $X=1715340 $Y=2015038
X220 6898 2 6869 6833 4 NAND2BX1 $T=1746360 2075920 1 180 $X=1743720 $Y=2075518
X221 7167 2 7208 7058 4 NAND2BX1 $T=1816980 2005360 1 180 $X=1814340 $Y=2004958
X222 7323 2 7328 7297 4 NAND2BX1 $T=1838100 2035600 0 180 $X=1835460 $Y=2030160
X223 7324 2 7329 7316 4 NAND2BX1 $T=1838100 2106160 0 180 $X=1835460 $Y=2100720
X224 7351 2 7354 7301 4 NAND2BX1 $T=1843380 2075920 0 180 $X=1840740 $Y=2070480
X225 7588 2 7566 7503 4 NAND2BX1 $T=1883640 2015440 1 180 $X=1881000 $Y=2015038
X226 7563 2 7603 7683 4 NAND2BX1 $T=1900800 2065840 1 0 $X=1900798 $Y=2060400
X227 7865 2 7864 7863 4 NAND2BX1 $T=1942380 2096080 1 180 $X=1939740 $Y=2095678
X228 7869 2 7877 7873 4 NAND2BX1 $T=1950300 1995280 0 0 $X=1950298 $Y=1994878
X229 7895 2 7907 7830 4 NAND2BX1 $T=1958220 2126320 1 0 $X=1958218 $Y=2120880
X230 8007 2 7984 7982 4 NAND2BX1 $T=1967460 2045680 0 180 $X=1964820 $Y=2040240
X231 554 2 8114 8116 4 NAND2BX1 $T=1994520 2217040 1 0 $X=1994518 $Y=2211600
X232 8114 2 554 8133 4 NAND2BX1 $T=1999140 2217040 0 0 $X=1999138 $Y=2216638
X233 8189 2 8190 8191 4 NAND2BX1 $T=2001120 2126320 0 0 $X=2001118 $Y=2125918
X234 8303 2 8281 8261 4 NAND2BX1 $T=2023560 2035600 1 180 $X=2020920 $Y=2035198
X235 8306 2 8290 8244 4 NAND2BX1 $T=2026200 2086000 0 180 $X=2023560 $Y=2080560
X236 8332 2 8312 8310 4 NAND2BX1 $T=2031480 2196880 0 180 $X=2028840 $Y=2191440
X237 577 2 576 8337 4 NAND2BX1 $T=2047320 1995280 0 180 $X=2044680 $Y=1989840
X238 8552 2 8555 8544 4 NAND2BX1 $T=2080980 2206960 0 0 $X=2080978 $Y=2206558
X239 8671 2 8609 8629 4 NAND2BX1 $T=2100780 2206960 0 180 $X=2098140 $Y=2201520
X240 8697 2 8691 8676 4 NAND2BX1 $T=2106060 2156560 1 180 $X=2103420 $Y=2156158
X241 8701 2 8724 8747 4 NAND2BX1 $T=2121900 2136400 1 180 $X=2119260 $Y=2135998
X242 8891 2 8876 8824 4 NAND2BX1 $T=2148960 2035600 0 180 $X=2146320 $Y=2030160
X243 8968 2 8972 8928 4 NAND2BX1 $T=2167440 2035600 0 180 $X=2164800 $Y=2030160
X244 9684 2 9683 9581 4 NAND2BX1 $T=2307360 2206960 1 180 $X=2304720 $Y=2206558
X245 10078 2 10139 10220 4 NAND2BX1 $T=2410980 2126320 1 0 $X=2410978 $Y=2120880
X246 10202 2 10199 10163 4 NAND2BX1 $T=2416920 2186800 1 180 $X=2414280 $Y=2186398
X247 693 2 10522 691 4 NAND2BX1 $T=2481600 1995280 0 180 $X=2478960 $Y=1989840
X248 10461 2 10440 10498 4 NAND2BX1 $T=2484240 2116240 0 180 $X=2481600 $Y=2110800
X249 707 2 713 10914 4 NAND2BX1 $T=2533740 2227120 1 0 $X=2533738 $Y=2221680
X250 74 73 2 69 4 779 OAI21X1 $T=766920 2227120 1 180 $X=763620 $Y=2226718
X251 2397 2445 2 2359 4 99 OAI21X1 $T=840180 2227120 0 180 $X=836880 $Y=2221680
X252 3110 3107 2 3059 4 3062 OAI21X1 $T=958980 2045680 1 0 $X=958978 $Y=2040240
X253 5077 5124 2 5019 4 5130 OAI21X1 $T=1360260 2146480 0 0 $X=1360258 $Y=2146078
X254 6054 6056 2 6059 4 5977 OAI21X1 $T=1563540 2065840 1 0 $X=1563538 $Y=2060400
X255 6710 6763 2 6743 4 6760 OAI21X1 $T=1718640 2045680 1 180 $X=1715340 $Y=2045278
X256 7059 7167 2 7208 4 7165 OAI21X1 $T=1807740 2005360 0 0 $X=1807738 $Y=2004958
X257 7502 7525 2 7523 4 7615 OAI21X1 $T=1885620 2045680 0 0 $X=1885618 $Y=2045278
X258 7865 7845 2 7864 4 7829 OAI21X1 $T=1941060 2106160 0 0 $X=1941058 $Y=2105758
X259 8303 8260 2 8281 4 8307 OAI21X1 $T=2026860 2035600 0 0 $X=2026858 $Y=2035198
X260 8552 8519 2 8555 4 8674 OAI21X1 $T=2082300 2217040 1 0 $X=2082298 $Y=2211600
X261 9603 9542 2 653 4 9662 OAI21X1 $T=2299440 1995280 1 0 $X=2299438 $Y=1989840
X262 10199 10335 2 10433 4 10390 OAI21X1 $T=2457840 2186800 0 0 $X=2457838 $Y=2186398
X263 728 724 2 720 4 725 OAI21X1 $T=2582580 1995280 1 180 $X=2579280 $Y=1994878
X264 2359 2 2353 2337 4 2354 OAI21XL $T=824340 2206960 1 180 $X=821700 $Y=2206558
X265 2684 2 2666 2667 4 2668 OAI21XL $T=887040 2146480 1 180 $X=884400 $Y=2146078
X266 2721 2 2717 2666 4 2713 OAI21XL $T=894960 2146480 1 180 $X=892320 $Y=2146078
X267 3327 2 3226 3159 4 3228 OAI21XL $T=991320 2035600 0 180 $X=988680 $Y=2030160
X268 3231 2 3260 3327 4 3254 OAI21XL $T=997260 2055760 0 180 $X=994620 $Y=2050320
X269 3364 2 3273 3433 4 3271 OAI21XL $T=998580 2186800 1 180 $X=995940 $Y=2186398
X270 3438 2 3409 3411 4 3229 OAI21XL $T=1016400 2055760 1 180 $X=1013760 $Y=2055358
X271 3488 2 3450 3494 4 3511 OAI21XL $T=1032240 2106160 0 0 $X=1032238 $Y=2105758
X272 3541 2 3538 3508 4 3466 OAI21XL $T=1044780 2005360 1 180 $X=1042140 $Y=2004958
X273 3565 2 3549 3640 4 3497 OAI21XL $T=1046760 2025520 0 180 $X=1044120 $Y=2020080
X274 3563 2 3538 3549 4 3548 OAI21XL $T=1048080 2015440 1 180 $X=1045440 $Y=2015038
X275 3494 2 3560 3566 4 3449 OAI21XL $T=1046100 2106160 1 0 $X=1046098 $Y=2100720
X276 3915 2 3737 3781 4 3868 OAI21XL $T=1122660 2065840 0 180 $X=1120020 $Y=2060400
X277 3936 2 3988 3915 4 3984 OAI21XL $T=1141140 2065840 1 0 $X=1141138 $Y=2060400
X278 4483 2 4382 4443 4 4110 OAI21XL $T=1237500 2015440 1 180 $X=1234860 $Y=2015038
X279 4547 2 4534 4543 4 4504 OAI21XL $T=1248060 2096080 1 180 $X=1245420 $Y=2095678
X280 4659 2 4534 4661 4 4660 OAI21XL $T=1269180 2096080 1 0 $X=1269178 $Y=2090640
X281 4849 2 4741 4811 4 4720 OAI21XL $T=1301520 2116240 0 180 $X=1298880 $Y=2110800
X282 4949 2 4973 4978 4 4965 OAI21XL $T=1334520 2086000 1 0 $X=1334518 $Y=2080560
X283 4848 2 5012 5016 4 5015 OAI21XL $T=1342440 2065840 1 0 $X=1342438 $Y=2060400
X284 5024 2 5028 5038 4 277 OAI21XL $T=1346400 1995280 0 0 $X=1346398 $Y=1994878
X285 5038 2 5078 5126 4 5084 OAI21XL $T=1360920 1995280 0 0 $X=1360918 $Y=1994878
X286 4196 2 349 5929 4 5871 OAI21XL $T=1537140 2196880 1 0 $X=1537138 $Y=2191440
X287 364 2 4469 6053 4 5954 OAI21XL $T=1561560 2166640 0 0 $X=1561558 $Y=2166238
X288 6254 2 6246 6249 4 6195 OAI21XL $T=1605120 2005360 1 180 $X=1602480 $Y=2004958
X289 423 2 6787 6759 4 6761 OAI21XL $T=1721280 2015440 0 0 $X=1721278 $Y=2015038
X290 6898 2 6828 6869 4 6925 OAI21XL $T=1754280 2075920 1 180 $X=1751640 $Y=2075518
X291 7068 2 7040 7059 4 7056 OAI21XL $T=1789260 2015440 0 180 $X=1786620 $Y=2010000
X292 7324 2 7314 7329 4 7365 OAI21XL $T=1843380 2106160 1 0 $X=1843378 $Y=2100720
X293 7869 2 521 7877 4 7955 OAI21XL $T=1943700 2005360 1 0 $X=1943698 $Y=1999920
X294 8001 2 8056 8057 4 8069 OAI21XL $T=1980000 2106160 0 0 $X=1979998 $Y=2105758
X295 8079 2 540 547 4 8206 OAI21XL $T=1985940 2005360 0 0 $X=1985938 $Y=2004958
X296 8187 2 8189 8190 4 8192 OAI21XL $T=2000460 2136400 0 0 $X=2000458 $Y=2135998
X297 8306 2 8243 8290 4 8292 OAI21XL $T=2030160 2086000 1 0 $X=2030158 $Y=2080560
X298 8208 2 8332 8312 4 8335 OAI21XL $T=2036760 2196880 0 180 $X=2034120 $Y=2191440
X299 8525 2 8514 8457 4 8511 OAI21XL $T=2074380 2146480 1 180 $X=2071740 $Y=2146078
X300 8457 2 8522 8493 4 8548 OAI21XL $T=2075700 2136400 1 0 $X=2075698 $Y=2130960
X301 8587 2 8569 8584 4 8572 OAI21XL $T=2091540 2136400 1 0 $X=2091538 $Y=2130960
X302 8671 2 8667 8609 4 8720 OAI21XL $T=2104740 2206960 1 0 $X=2104738 $Y=2201520
X303 8697 2 8673 8691 4 8745 OAI21XL $T=2111340 2156560 0 0 $X=2111338 $Y=2156158
X304 8691 2 8701 8724 4 8694 OAI21XL $T=2113980 2136400 1 180 $X=2111340 $Y=2135998
X305 610 2 609 606 4 8849 OAI21XL $T=2136420 1995280 0 0 $X=2136418 $Y=1994878
X306 8882 2 8717 8926 4 9015 OAI21XL $T=2152920 2146480 1 0 $X=2152918 $Y=2141040
X307 9036 2 9025 9018 4 9082 OAI21XL $T=2178660 2156560 0 0 $X=2178658 $Y=2156158
X308 9540 2 9686 9531 4 9689 OAI21XL $T=2307360 2156560 0 0 $X=2307358 $Y=2156158
X309 9531 2 9698 9700 4 9733 OAI21XL $T=2327160 2146480 0 0 $X=2327158 $Y=2146078
X310 9879 2 9939 9938 4 10140 OAI21XL $T=2359500 2126320 0 0 $X=2359498 $Y=2125918
X311 10136 2 10078 10139 4 10184 OAI21XL $T=2403060 2126320 0 0 $X=2403058 $Y=2125918
X312 10298 2 10320 10322 4 10412 OAI21XL $T=2443320 2136400 1 0 $X=2443318 $Y=2130960
X313 10556 2 10442 10562 4 10500 OAI21XL $T=2486880 2126320 1 0 $X=2486878 $Y=2120880
X314 10440 2 10568 10570 4 10655 OAI21XL $T=2489520 2106160 1 0 $X=2489518 $Y=2100720
X315 10461 2 10325 10440 4 10569 OAI21XL $T=2492820 2116240 0 180 $X=2490180 $Y=2110800
X316 10322 2 10683 10684 4 10727 OAI21XL $T=2509980 2116240 0 0 $X=2509978 $Y=2115838
X317 704 2 10658 10726 4 705 OAI21XL $T=2513940 1995280 0 0 $X=2513938 $Y=1994878
X318 10610 2 10442 10656 4 10722 OAI21XL $T=2520540 2126320 0 0 $X=2520538 $Y=2125918
X319 707 2 711 713 4 10790 OAI21XL $T=2530440 2227120 0 0 $X=2530438 $Y=2226718
X320 10746 2 10442 10911 4 10847 OAI21XL $T=2541660 2116240 0 0 $X=2541658 $Y=2115838
X321 10982 2 10442 10990 4 10880 OAI21XL $T=2554860 2126320 0 180 $X=2552220 $Y=2120880
X322 10941 2 10972 10981 4 10984 OAI21XL $T=2553540 2096080 0 0 $X=2553538 $Y=2095678
X323 11022 2 10442 11026 4 11001 OAI21XL $T=2560140 2116240 1 180 $X=2557500 $Y=2115838
X324 11043 2 10442 11095 4 11060 OAI21XL $T=2579280 2126320 1 0 $X=2579278 $Y=2120880
X325 10987 2 11094 11004 4 11110 OAI21XL $T=2579940 2086000 1 0 $X=2579938 $Y=2080560
X326 11133 2 10442 11129 4 11160 OAI21XL $T=2588520 2116240 0 0 $X=2588518 $Y=2115838
X327 2519 2445 780 2 4 XOR2X4 $T=851400 2227120 0 0 $X=851398 $Y=2226718
X328 2616 2655 105 2 4 XOR2X4 $T=875160 2196880 1 0 $X=875158 $Y=2191440
X329 5108 5099 5152 2 4 XOR2X4 $T=1358280 2196880 0 0 $X=1358278 $Y=2196478
X330 7613 7589 496 2 4 XOR2X4 $T=1896180 2096080 1 180 $X=1884960 $Y=2095678
X331 7779 7812 518 2 4 XOR2X4 $T=1922580 2166640 1 0 $X=1922578 $Y=2161200
X332 7828 7851 529 2 4 XOR2X4 $T=1933800 2186800 1 0 $X=1933798 $Y=2181360
X333 7863 7845 515 2 4 XOR2X4 $T=1945680 2096080 0 180 $X=1934460 $Y=2090640
X334 8070 551 552 2 4 XOR2X4 $T=1983300 2217040 0 0 $X=1983298 $Y=2216638
X335 557 531 560 2 4 XOR2X4 $T=1997160 2227120 0 0 $X=1997158 $Y=2226718
X336 9510 9429 646 2 4 XOR2X4 $T=2277660 2206960 0 180 $X=2266440 $Y=2201520
X337 9655 9581 652 2 4 XOR2X4 $T=2300760 2206960 0 180 $X=2289540 $Y=2201520
X338 9914 9910 665 2 4 XOR2X4 $T=2358840 2196880 0 180 $X=2347620 $Y=2191440
X339 9994 9971 671 2 4 XOR2X4 $T=2374680 2196880 0 180 $X=2363460 $Y=2191440
X340 10163 10141 679 2 4 XOR2X4 $T=2409000 2186800 0 180 $X=2397780 $Y=2181360
X341 690 686 10415 2 4 XOR2X4 $T=2467080 2227120 0 180 $X=2455860 $Y=2221680
X342 694 692 10523 2 4 XOR2X4 $T=2490840 2227120 0 180 $X=2479620 $Y=2221680
X343 695 698 10685 2 4 XOR2X4 $T=2499420 2227120 1 0 $X=2499418 $Y=2221680
X344 2636 2 4 2659 INVX1 $T=878460 2136400 1 0 $X=878458 $Y=2130960
X345 2708 2 4 2679 INVX1 $T=891660 2116240 0 0 $X=891658 $Y=2115838
X346 2679 2 4 2751 INVX1 $T=899580 2126320 0 0 $X=899578 $Y=2125918
X347 2716 2 4 2790 INVX1 $T=904860 2126320 1 0 $X=904858 $Y=2120880
X348 2788 2 4 2829 INVX1 $T=906180 2005360 1 0 $X=906178 $Y=1999920
X349 2826 2 4 2834 INVX1 $T=918720 2005360 1 180 $X=917400 $Y=2004958
X350 2844 2 4 2845 INVX1 $T=918720 2086000 1 180 $X=917400 $Y=2085598
X351 2839 2 4 2883 INVX1 $T=918060 2106160 1 0 $X=918058 $Y=2100720
X352 2928 2 4 2888 INVX1 $T=935220 2096080 1 180 $X=933900 $Y=2095678
X353 2956 2 4 2984 INVX1 $T=939180 2176720 0 0 $X=939178 $Y=2176318
X354 3058 2 4 3081 INVX1 $T=949080 2196880 1 0 $X=949078 $Y=2191440
X355 3066 2 4 3061 INVX1 $T=955680 2025520 1 180 $X=954360 $Y=2025118
X356 3118 2 4 3109 INVX1 $T=960960 2186800 1 180 $X=959640 $Y=2186398
X357 3145 2 4 3119 INVX1 $T=964920 2126320 0 180 $X=963600 $Y=2120880
X358 3084 2 4 3085 INVX1 $T=964920 2176720 1 0 $X=964918 $Y=2171280
X359 116 2 4 3063 INVX1 $T=966240 2217040 1 180 $X=964920 $Y=2216638
X360 3144 2 4 3158 INVX1 $T=970200 2065840 0 0 $X=970198 $Y=2065438
X361 67 2 4 118 INVX1 $T=978120 2005360 1 0 $X=978118 $Y=1999920
X362 3195 2 4 3136 INVX1 $T=981420 2126320 1 180 $X=980100 $Y=2125918
X363 3200 2 4 3218 INVX1 $T=982740 2065840 0 0 $X=982738 $Y=2065438
X364 3274 2 4 3278 INVX1 $T=997920 2196880 1 180 $X=996600 $Y=2196478
X365 3363 2 4 3366 INVX1 $T=1007160 2126320 1 0 $X=1007158 $Y=2120880
X366 3409 2 4 3435 INVX1 $T=1017060 2065840 1 0 $X=1017058 $Y=2060400
X367 3450 2 4 3442 INVX1 $T=1026300 2106160 0 180 $X=1024980 $Y=2100720
X368 3461 2 4 3513 INVX1 $T=1032240 2005360 1 0 $X=1032238 $Y=1999920
X369 3443 2 4 3431 INVX1 $T=1034220 2116240 0 180 $X=1032900 $Y=2110800
X370 3482 2 4 3469 INVX1 $T=1036860 2176720 1 180 $X=1035540 $Y=2176318
X371 3519 2 4 3543 INVX1 $T=1038180 2156560 0 0 $X=1038178 $Y=2156158
X372 3438 2 4 3535 INVX1 $T=1039500 2055760 0 0 $X=1039498 $Y=2055358
X373 3500 2 4 3538 INVX1 $T=1040820 2015440 0 0 $X=1040818 $Y=2015038
X374 3483 2 4 3619 INVX1 $T=1048740 2186800 1 0 $X=1048738 $Y=2181360
X375 3618 2 4 3514 INVX1 $T=1050060 2116240 1 180 $X=1048740 $Y=2115838
X376 3464 2 4 3659 INVX1 $T=1061940 2065840 0 0 $X=1061938 $Y=2065438
X377 3658 2 4 3703 INVX1 $T=1067220 2075920 1 0 $X=1067218 $Y=2070480
X378 125 2 4 137 INVX1 $T=1074480 2015440 1 0 $X=1074478 $Y=2010000
X379 3758 2 4 3739 INVX1 $T=1087020 2035600 0 180 $X=1085700 $Y=2030160
X380 3787 2 4 3725 INVX1 $T=1092960 2035600 0 0 $X=1092958 $Y=2035198
X381 3815 2 4 128 INVX1 $T=1101540 2075920 0 180 $X=1100220 $Y=2070480
X382 3861 2 4 3780 INVX1 $T=1108800 2035600 1 0 $X=1108798 $Y=2030160
X383 3737 2 4 3880 INVX1 $T=1111440 2075920 1 0 $X=1111438 $Y=2070480
X384 3917 2 4 3919 INVX1 $T=1123980 2015440 0 0 $X=1123978 $Y=2015038
X385 3666 2 4 3765 INVX1 $T=1152360 2096080 0 180 $X=1151040 $Y=2090640
X386 3818 2 4 3696 INVX1 $T=1153020 2126320 0 180 $X=1151700 $Y=2120880
X387 3988 2 4 3879 INVX1 $T=1158300 2065840 1 0 $X=1158298 $Y=2060400
X388 4110 2 4 3988 INVX1 $T=1162260 2055760 0 180 $X=1160940 $Y=2050320
X389 149 2 4 3638 INVX1 $T=1194600 2136400 1 0 $X=1194598 $Y=2130960
X390 132 2 4 4604 INVX1 $T=1252680 2035600 0 0 $X=1252678 $Y=2035198
X391 4507 2 4 4605 INVX1 $T=1252680 2086000 1 0 $X=1252678 $Y=2080560
X392 4547 2 4 4535 INVX1 $T=1255320 2106160 0 0 $X=1255318 $Y=2105758
X393 4720 2 4 4534 INVX1 $T=1269840 2106160 0 180 $X=1268520 $Y=2100720
X394 248 2 4 246 INVX1 $T=1280400 1995280 0 180 $X=1279080 $Y=1989840
X395 4735 2 4 4721 INVX1 $T=1287000 2126320 1 0 $X=1286998 $Y=2120880
X396 4741 2 4 4702 INVX1 $T=1288320 2116240 1 180 $X=1287000 $Y=2115838
X397 4786 2 4 4752 INVX1 $T=1296900 2015440 1 180 $X=1295580 $Y=2015038
X398 4797 2 4 4794 INVX1 $T=1300860 2126320 1 180 $X=1299540 $Y=2125918
X399 4848 2 4 4888 INVX1 $T=1319340 2075920 0 180 $X=1318020 $Y=2070480
X400 252 2 4 255 INVX1 $T=1323300 2015440 1 0 $X=1323298 $Y=2010000
X401 4891 2 4 4976 INVX1 $T=1323300 2217040 1 0 $X=1323298 $Y=2211600
X402 4913 2 4 4956 INVX1 $T=1332540 2146480 1 180 $X=1331220 $Y=2146078
X403 4995 2 4 5000 INVX1 $T=1339140 2196880 0 0 $X=1339138 $Y=2196478
X404 5015 2 4 5028 INVX1 $T=1344420 1995280 1 180 $X=1343100 $Y=1994878
X405 4994 2 4 5027 INVX1 $T=1347060 2196880 1 0 $X=1347058 $Y=2191440
X406 5085 2 4 5124 INVX1 $T=1364220 2116240 0 180 $X=1362900 $Y=2110800
X407 285 2 4 4320 INVX1 $T=1368840 2096080 0 180 $X=1367520 $Y=2090640
X408 262 2 4 268 INVX1 $T=1386000 2176720 0 0 $X=1385998 $Y=2176318
X409 5230 2 4 5234 INVX1 $T=1391940 2106160 1 0 $X=1391938 $Y=2100720
X410 5343 2 4 5404 INVX1 $T=1415040 2075920 1 0 $X=1415038 $Y=2070480
X411 218 2 4 5209 INVX1 $T=1445400 2086000 0 180 $X=1444080 $Y=2080560
X412 309 2 4 5598 INVX1 $T=1457940 2035600 1 0 $X=1457938 $Y=2030160
X413 5871 2 4 5920 INVX1 $T=1524600 2217040 0 0 $X=1524598 $Y=2216638
X414 218 2 4 5953 INVX1 $T=1542420 2086000 1 0 $X=1542418 $Y=2080560
X415 5982 2 4 5981 INVX1 $T=1551000 2096080 0 0 $X=1550998 $Y=2095678
X416 310 2 4 346 INVX1 $T=1552980 2055760 1 0 $X=1552978 $Y=2050320
X417 363 2 4 5508 INVX1 $T=1582020 2106160 1 0 $X=1582018 $Y=2100720
X418 325 2 4 297 INVX1 $T=1598520 2015440 1 180 $X=1597200 $Y=2015038
X419 6257 2 4 6189 INVX1 $T=1604460 2045680 0 180 $X=1603140 $Y=2040240
X420 373 2 4 6216 INVX1 $T=1611720 2116240 1 180 $X=1610400 $Y=2115838
X421 6297 2 4 380 INVX1 $T=1614360 2217040 1 180 $X=1613040 $Y=2216638
X422 383 2 4 6287 INVX1 $T=1615020 2075920 0 180 $X=1613700 $Y=2070480
X423 6335 2 4 6324 INVX1 $T=1622280 2015440 0 180 $X=1620960 $Y=2010000
X424 6405 2 4 370 INVX1 $T=1640760 2156560 1 180 $X=1639440 $Y=2156158
X425 6481 2 4 6334 INVX1 $T=1641420 2015440 1 180 $X=1640100 $Y=2015038
X426 310 2 4 389 INVX1 $T=1644720 2227120 1 0 $X=1644718 $Y=2221680
X427 400 2 4 343 INVX1 $T=1659240 2217040 0 180 $X=1657920 $Y=2211600
X428 6697 2 4 6709 INVX1 $T=1702800 2005360 0 0 $X=1702798 $Y=2004958
X429 6715 2 4 6771 INVX1 $T=1716000 2075920 1 0 $X=1715998 $Y=2070480
X430 310 2 4 437 INVX1 $T=1728540 2217040 0 0 $X=1728538 $Y=2216638
X431 325 2 4 430 INVX1 $T=1734480 2227120 0 180 $X=1733160 $Y=2221680
X432 227 2 4 314 INVX1 $T=1735140 1995280 1 0 $X=1735138 $Y=1989840
X433 6850 2 4 6853 INVX1 $T=1741740 2055760 0 0 $X=1741738 $Y=2055358
X434 349 2 4 440 INVX1 $T=1745040 2106160 1 0 $X=1745038 $Y=2100720
X435 6986 2 4 6991 INVX1 $T=1776060 2096080 0 0 $X=1776058 $Y=2095678
X436 7046 2 4 7091 INVX1 $T=1783980 2086000 0 0 $X=1783978 $Y=2085598
X437 7047 2 4 7053 INVX1 $T=1793880 2055760 0 0 $X=1793878 $Y=2055358
X438 7166 2 4 7216 INVX1 $T=1815000 2116240 0 0 $X=1814998 $Y=2115838
X439 7257 2 4 7211 INVX1 $T=1821600 2096080 0 180 $X=1820280 $Y=2090640
X440 7260 2 4 7296 INVX1 $T=1830840 2025520 1 0 $X=1830838 $Y=2020080
X441 7297 2 4 7300 INVX1 $T=1830840 2035600 0 0 $X=1830838 $Y=2035198
X442 7219 2 4 7314 INVX1 $T=1830840 2106160 1 0 $X=1830838 $Y=2100720
X443 7454 2 4 7430 INVX1 $T=1860540 2005360 1 180 $X=1859220 $Y=2004958
X444 7592 2 4 7616 INVX1 $T=1890900 2116240 1 0 $X=1890898 $Y=2110800
X445 499 2 4 7705 INVX1 $T=1894860 2217040 0 0 $X=1894858 $Y=2216638
X446 7635 2 4 7688 INVX1 $T=1901460 2086000 0 0 $X=1901458 $Y=2085598
X447 7690 2 4 7686 INVX1 $T=1904760 2106160 0 180 $X=1903440 $Y=2100720
X448 509 2 4 7730 INVX1 $T=1915320 2217040 0 180 $X=1914000 $Y=2211600
X449 7755 2 4 7772 INVX1 $T=1917960 2045680 0 180 $X=1916640 $Y=2040240
X450 519 2 4 7802 INVX1 $T=1933800 2206960 0 180 $X=1932480 $Y=2201520
X451 7788 2 4 7846 INVX1 $T=1935120 2055760 1 0 $X=1935118 $Y=2050320
X452 512 2 4 7872 INVX1 $T=1940400 2206960 0 0 $X=1940398 $Y=2206558
X453 7955 2 4 8001 INVX1 $T=1957560 2075920 0 0 $X=1957558 $Y=2075518
X454 7962 2 4 7961 INVX1 $T=1958880 2045680 1 0 $X=1958878 $Y=2040240
X455 8025 2 4 8024 INVX1 $T=1973400 2096080 0 0 $X=1973398 $Y=2095678
X456 8069 2 4 8187 INVX1 $T=1984620 2116240 1 0 $X=1984618 $Y=2110800
X457 8188 2 4 8209 INVX1 $T=2000460 2176720 0 0 $X=2000458 $Y=2176318
X458 556 2 4 8112 INVX1 $T=2001120 2227120 1 0 $X=2001118 $Y=2221680
X459 8234 2 4 8215 INVX1 $T=2011020 2106160 1 0 $X=2011018 $Y=2100720
X460 8258 2 4 8239 INVX1 $T=2017620 2015440 1 180 $X=2016300 $Y=2015038
X461 8278 2 4 8263 INVX1 $T=2020260 2156560 1 180 $X=2018940 $Y=2156158
X462 8305 2 4 8322 INVX1 $T=2026860 2126320 1 0 $X=2026858 $Y=2120880
X463 8327 2 4 8329 INVX1 $T=2032140 2156560 1 0 $X=2032138 $Y=2151120
X464 8398 2 4 8405 INVX1 $T=2047980 2186800 1 0 $X=2047978 $Y=2181360
X465 8439 2 4 8473 INVX1 $T=2063820 2206960 0 0 $X=2063818 $Y=2206558
X466 8515 2 4 8516 INVX1 $T=2073720 2176720 1 0 $X=2073718 $Y=2171280
X467 587 2 4 8546 INVX1 $T=2076360 2015440 0 0 $X=2076358 $Y=2015038
X468 590 2 4 8588 INVX1 $T=2084280 1995280 0 0 $X=2084278 $Y=1994878
X469 8572 2 4 8673 INVX1 $T=2086920 2156560 0 0 $X=2086918 $Y=2156158
X470 8595 2 4 8608 INVX1 $T=2092200 2186800 0 0 $X=2092198 $Y=2186398
X471 8674 2 4 8667 INVX1 $T=2102760 2206960 0 0 $X=2102758 $Y=2206558
X472 8695 2 4 781 INVX1 $T=2106720 2227120 1 180 $X=2105400 $Y=2226718
X473 8740 2 4 8703 INVX1 $T=2125200 2015440 0 180 $X=2123880 $Y=2010000
X474 8717 2 4 8803 INVX1 $T=2127840 2146480 1 0 $X=2127838 $Y=2141040
X475 8784 2 4 607 INVX1 $T=2129160 2196880 1 0 $X=2129158 $Y=2191440
X476 8823 2 4 8827 INVX1 $T=2137080 2146480 0 0 $X=2137078 $Y=2146078
X477 8851 2 4 613 INVX1 $T=2143020 2196880 1 0 $X=2143018 $Y=2191440
X478 8890 2 4 8930 INVX1 $T=2149620 2156560 1 0 $X=2149618 $Y=2151120
X479 8891 2 4 8925 INVX1 $T=2156880 2035600 0 180 $X=2155560 $Y=2030160
X480 8975 2 4 8987 INVX1 $T=2172720 2206960 0 0 $X=2172718 $Y=2206558
X481 9015 2 4 9025 INVX1 $T=2173380 2146480 0 0 $X=2173378 $Y=2146078
X482 9011 2 4 8989 INVX1 $T=2173380 2186800 1 0 $X=2173378 $Y=2181360
X483 9037 2 4 9024 INVX1 $T=2179980 2196880 1 180 $X=2178660 $Y=2196478
X484 9108 2 4 9064 INVX1 $T=2193180 2176720 1 180 $X=2191860 $Y=2176318
X485 9190 2 4 9168 INVX1 $T=2209020 2196880 0 180 $X=2207700 $Y=2191440
X486 9181 2 4 9255 INVX1 $T=2217600 2025520 1 0 $X=2217598 $Y=2020080
X487 9169 2 4 9249 INVX1 $T=2218920 2227120 1 0 $X=2218918 $Y=2221680
X488 9269 2 4 9278 INVX1 $T=2225520 2025520 1 0 $X=2225518 $Y=2020080
X489 9319 2 4 9333 INVX1 $T=2238720 2166640 1 0 $X=2238718 $Y=2161200
X490 9316 2 4 9322 INVX1 $T=2238720 2186800 0 0 $X=2238718 $Y=2186398
X491 9281 2 4 9338 INVX1 $T=2242020 2146480 0 0 $X=2242018 $Y=2146078
X492 9342 2 4 9405 INVX1 $T=2246640 2206960 1 0 $X=2246638 $Y=2201520
X493 9331 2 4 9404 INVX1 $T=2251920 2156560 1 180 $X=2250600 $Y=2156158
X494 9425 2 4 9453 INVX1 $T=2259840 2025520 1 0 $X=2259838 $Y=2020080
X495 9488 2 4 9431 INVX1 $T=2267760 2217040 1 180 $X=2266440 $Y=2216638
X496 9337 2 4 9494 INVX1 $T=2273040 2146480 1 0 $X=2273038 $Y=2141040
X497 9522 2 4 9489 INVX1 $T=2280300 2186800 0 0 $X=2280298 $Y=2186398
X498 9498 2 4 9686 INVX1 $T=2310660 2156560 0 180 $X=2309340 $Y=2151120
X499 658 2 4 9666 INVX1 $T=2315940 2005360 1 180 $X=2314620 $Y=2004958
X500 9725 2 4 9734 INVX1 $T=2317260 1995280 0 0 $X=2317258 $Y=1994878
X501 9775 2 4 9699 INVX1 $T=2327820 2206960 0 180 $X=2326500 $Y=2201520
X502 9878 2 4 9859 INVX1 $T=2347620 2176720 1 180 $X=2346300 $Y=2176318
X503 9916 2 4 9918 INVX1 $T=2354880 2176720 1 0 $X=2354878 $Y=2171280
X504 9930 2 4 9957 INVX1 $T=2357520 2206960 1 0 $X=2357518 $Y=2201520
X505 10018 2 4 10012 INVX1 $T=2382600 2217040 0 0 $X=2382598 $Y=2216638
X506 10015 2 4 10141 INVX1 $T=2405700 2186800 0 0 $X=2405698 $Y=2186398
X507 10246 2 4 10232 INVX1 $T=2425500 2176720 0 180 $X=2424180 $Y=2171280
X508 10202 2 4 10276 INVX1 $T=2434740 2186800 0 0 $X=2434738 $Y=2186398
X509 10222 2 4 10294 INVX1 $T=2437380 2126320 0 0 $X=2437378 $Y=2125918
X510 10317 2 4 10297 INVX1 $T=2444640 2186800 1 180 $X=2443320 $Y=2186398
X511 10411 2 4 10414 INVX1 $T=2455860 2035600 0 0 $X=2455858 $Y=2035198
X512 10230 2 4 10486 INVX1 $T=2463780 2136400 0 0 $X=2463778 $Y=2135998
X513 10470 2 4 10472 INVX1 $T=2469060 2045680 0 0 $X=2469058 $Y=2045278
X514 10486 2 4 10542 INVX1 $T=2476320 2136400 1 0 $X=2476318 $Y=2130960
X515 10540 2 4 10462 INVX1 $T=2486220 2176720 1 180 $X=2484900 $Y=2176318
X516 10325 2 4 10608 INVX1 $T=2492160 2116240 0 0 $X=2492158 $Y=2115838
X517 10298 2 4 10560 INVX1 $T=2504040 2136400 1 180 $X=2502720 $Y=2135998
X518 10681 2 4 10682 INVX1 $T=2508000 2055760 1 0 $X=2507998 $Y=2050320
X519 10322 2 4 10657 INVX1 $T=2510640 2136400 1 0 $X=2510638 $Y=2130960
X520 10815 2 4 10662 INVX1 $T=2517240 2025520 0 180 $X=2515920 $Y=2020080
X521 708 2 4 10886 INVX1 $T=2537040 2227120 0 0 $X=2537038 $Y=2226718
X522 10782 2 4 10746 INVX1 $T=2543640 2116240 0 180 $X=2542320 $Y=2110800
X523 711 2 4 10917 INVX1 $T=2544960 2227120 0 0 $X=2544958 $Y=2226718
X524 10727 2 4 10911 INVX1 $T=2548920 2116240 1 180 $X=2547600 $Y=2115838
X525 10922 2 4 10989 INVX1 $T=2555520 1995280 1 0 $X=2555518 $Y=1989840
X526 10980 2 4 10973 INVX1 $T=2562780 2065840 0 0 $X=2562778 $Y=2065438
X527 10941 2 4 11029 INVX1 $T=2562780 2106160 1 0 $X=2562778 $Y=2100720
X528 11021 2 4 11064 INVX1 $T=2573340 2035600 0 0 $X=2573338 $Y=2035198
X529 11090 2 4 11092 INVX1 $T=2578620 2035600 0 0 $X=2578618 $Y=2035198
X530 11065 2 4 11155 INVX1 $T=2597100 2096080 1 0 $X=2597098 $Y=2090640
X531 11163 2 4 11227 INVX1 $T=2599740 2045680 0 0 $X=2599738 $Y=2045278
X532 11226 2 4 736 INVX1 $T=2609640 1995280 1 0 $X=2609638 $Y=1989840
X533 11154 2 4 11290 INVX1 $T=2612940 2005360 1 0 $X=2612938 $Y=1999920
X534 2384 2451 4 2354 2444 2 AOI21X2 $T=846120 2206960 1 180 $X=841500 $Y=2206558
X535 2831 2685 4 2668 2632 2 AOI21X2 $T=889680 2176720 0 180 $X=885060 $Y=2171280
X536 3085 3139 4 3081 3111 2 AOI21X2 $T=966900 2196880 0 180 $X=962280 $Y=2191440
X537 3199 3229 4 3228 3237 2 AOI21X2 $T=988020 2065840 1 0 $X=988018 $Y=2060400
X538 3500 3510 4 3497 3450 2 AOI21X2 $T=1037520 2035600 0 180 $X=1032900 $Y=2030160
X539 3898 3879 4 3868 3532 2 AOI21X2 $T=1113420 2065840 0 180 $X=1108800 $Y=2060400
X540 5000 4908 4 4976 4992 2 AOI21X2 $T=1341120 2217040 0 180 $X=1336500 $Y=2211600
X541 5961 5977 4 5981 5930 2 AOI21X2 $T=1547700 2086000 1 0 $X=1547698 $Y=2080560
X542 6764 6760 4 6853 6866 2 AOI21X2 $T=1739100 2055760 1 0 $X=1739098 $Y=2050320
X543 7021 7045 4 7053 7069 2 AOI21X2 $T=1783320 2055760 0 0 $X=1783318 $Y=2055358
X544 7170 7211 4 7216 7187 2 AOI21X2 $T=1811040 2106160 0 0 $X=1811038 $Y=2105758
X545 7686 7607 4 7616 7681 2 AOI21X2 $T=1900140 2116240 0 180 $X=1895520 $Y=2110800
X546 7614 7730 4 7705 7727 2 AOI21X2 $T=1913340 2217040 1 180 $X=1908720 $Y=2216638
X547 7810 7777 4 7846 7878 2 AOI21X2 $T=1945020 2055760 0 180 $X=1940400 $Y=2050320
X548 7962 8023 4 8028 8005 2 AOI21X2 $T=1971420 2045680 1 0 $X=1971418 $Y=2040240
X549 551 553 4 8112 8114 2 AOI21X2 $T=1992540 2227120 1 0 $X=1992538 $Y=2221680
X550 615 8970 4 8987 8992 2 AOI21X2 $T=2170080 2206960 0 180 $X=2165460 $Y=2201520
X551 9421 9344 4 9405 9429 2 AOI21X2 $T=2258520 2206960 0 180 $X=2253900 $Y=2201520
X552 9422 9405 4 9431 9457 2 AOI21X2 $T=2256540 2217040 0 0 $X=2256538 $Y=2216638
X553 9910 9917 4 9957 9971 2 AOI21X2 $T=2364120 2206960 1 0 $X=2364118 $Y=2201520
X554 672 9957 4 10012 10011 2 AOI21X2 $T=2374680 2217040 1 0 $X=2374678 $Y=2211600
X555 4 2097 2093 77 2 NOR2X1 $T=767580 2196880 1 0 $X=767578 $Y=2191440
X556 4 2565 2560 2557 2 NOR2X1 $T=861300 2146480 1 180 $X=859320 $Y=2146078
X557 4 2588 2422 2540 2 NOR2X1 $T=867240 2176720 0 180 $X=865260 $Y=2171280
X558 4 2603 2630 2684 2 NOR2X1 $T=876480 2156560 1 0 $X=876478 $Y=2151120
X559 4 2721 2684 2685 2 NOR2X1 $T=888360 2156560 1 180 $X=886380 $Y=2156158
X560 4 2828 2786 2788 2 NOR2X1 $T=915420 2005360 0 180 $X=913440 $Y=1999920
X561 4 108 2892 2868 2 NOR2X1 $T=927300 2227120 0 180 $X=925320 $Y=2221680
X562 4 93 2885 2976 2 NOR2X1 $T=934560 1995280 0 0 $X=934558 $Y=1994878
X563 4 2421 55 3107 2 NOR2X1 $T=950400 2045680 0 0 $X=950398 $Y=2045278
X564 4 3088 2804 3084 2 NOR2X1 $T=958980 2146480 0 0 $X=958978 $Y=2146078
X565 4 3145 3166 3184 2 NOR2X1 $T=973500 2146480 0 0 $X=973498 $Y=2146078
X566 4 3230 2977 3166 2 NOR2X1 $T=988680 2106160 1 0 $X=988678 $Y=2100720
X567 4 3409 3389 3186 2 NOR2X1 $T=1013760 2065840 0 180 $X=1011780 $Y=2060400
X568 4 3416 3122 3409 2 NOR2X1 $T=1017720 2045680 0 180 $X=1015740 $Y=2040240
X569 4 3481 3255 3389 2 NOR2X1 $T=1030920 2055760 1 0 $X=1030918 $Y=2050320
X570 4 3488 3560 3471 2 NOR2X1 $T=1047420 2116240 0 180 $X=1045440 $Y=2110800
X571 4 3565 3563 3510 2 NOR2X1 $T=1048080 2035600 0 180 $X=1046100 $Y=2030160
X572 4 3569 3564 3488 2 NOR2X1 $T=1048080 2086000 1 180 $X=1046100 $Y=2085598
X573 4 125 124 3541 2 NOR2X1 $T=1048080 1995280 0 0 $X=1048078 $Y=1994878
X574 4 3698 3626 3560 2 NOR2X1 $T=1056000 2106160 0 180 $X=1054020 $Y=2100720
X575 4 131 128 3486 2 NOR2X1 $T=1065900 1995280 1 180 $X=1063920 $Y=1994878
X576 4 3746 3681 3443 2 NOR2X1 $T=1071180 2116240 1 180 $X=1069200 $Y=2115838
X577 4 3725 3722 3683 2 NOR2X1 $T=1080420 2045680 0 180 $X=1078440 $Y=2040240
X578 4 3794 163 162 2 NOR2X1 $T=1110780 1995280 1 180 $X=1108800 $Y=1994878
X579 4 3737 3936 3898 2 NOR2X1 $T=1127940 2065840 1 0 $X=1127938 $Y=2060400
X580 4 3956 95 3936 2 NOR2X1 $T=1133220 2055760 1 0 $X=1133218 $Y=2050320
X581 4 140 3958 3935 2 NOR2X1 $T=1134540 2025520 1 0 $X=1134538 $Y=2020080
X582 4 139 3987 3959 2 NOR2X1 $T=1140480 2035600 0 0 $X=1140478 $Y=2035198
X583 4 208 207 211 2 NOR2X1 $T=1214400 2227120 1 0 $X=1214398 $Y=2221680
X584 4 4321 203 4382 2 NOR2X1 $T=1215060 2015440 0 0 $X=1215058 $Y=2015038
X585 4 4486 4480 228 2 NOR2X1 $T=1239480 2227120 1 0 $X=1239478 $Y=2221680
X586 4 231 233 4547 2 NOR2X1 $T=1250700 2116240 1 0 $X=1250698 $Y=2110800
X587 4 4605 4618 4661 2 NOR2X1 $T=1255320 2086000 0 0 $X=1255318 $Y=2085598
X588 4 247 238 236 2 NOR2X1 $T=1265880 1995280 1 180 $X=1263900 $Y=1994878
X589 4 4638 4541 245 2 NOR2X1 $T=1267860 2227120 1 0 $X=1267858 $Y=2221680
X590 4 4703 4683 4719 2 NOR2X1 $T=1279740 2096080 1 0 $X=1279738 $Y=2090640
X591 4 4719 4659 4730 2 NOR2X1 $T=1282380 2106160 1 0 $X=1282378 $Y=2100720
X592 4 252 262 4786 2 NOR2X1 $T=1313400 2025520 0 180 $X=1311420 $Y=2020080
X593 4 4851 4968 4970 2 NOR2X1 $T=1333200 2106160 0 0 $X=1333198 $Y=2105758
X594 4 4970 4973 4954 2 NOR2X1 $T=1335180 2096080 0 180 $X=1333200 $Y=2090640
X595 4 4980 4996 5024 2 NOR2X1 $T=1338480 2005360 1 0 $X=1338478 $Y=1999920
X596 4 3337 275 5077 2 NOR2X1 $T=1349040 2156560 0 0 $X=1349038 $Y=2156158
X597 4 5003 5074 4973 2 NOR2X1 $T=1352340 2096080 1 180 $X=1350360 $Y=2095678
X598 4 5024 5078 5081 2 NOR2X1 $T=1351680 2005360 1 0 $X=1351678 $Y=1999920
X599 4 5096 5123 5078 2 NOR2X1 $T=1361580 2005360 1 180 $X=1359600 $Y=2004958
X600 4 3702 345 5874 2 NOR2X1 $T=1517340 2075920 1 0 $X=1517338 $Y=2070480
X601 4 6058 4108 6054 2 NOR2X1 $T=1566840 2065840 1 180 $X=1564860 $Y=2065438
X602 4 6270 4637 6246 2 NOR2X1 $T=1603800 2015440 0 180 $X=1601820 $Y=2010000
X603 4 6770 424 6763 2 NOR2X1 $T=1719960 2035600 0 180 $X=1717980 $Y=2030160
X604 4 6807 6080 6787 2 NOR2X1 $T=1726560 2025520 1 180 $X=1724580 $Y=2025118
X605 4 6944 5741 6898 2 NOR2X1 $T=1758900 2075920 1 0 $X=1758898 $Y=2070480
X606 4 7026 457 6987 2 NOR2X1 $T=1783320 2035600 0 0 $X=1783318 $Y=2035198
X607 4 7068 7167 7163 2 NOR2X1 $T=1803780 2015440 0 180 $X=1801800 $Y=2010000
X608 4 7189 470 7068 2 NOR2X1 $T=1803780 2015440 1 180 $X=1801800 $Y=2015038
X609 4 7168 469 7090 2 NOR2X1 $T=1803120 2045680 1 0 $X=1803118 $Y=2040240
X610 4 8024 541 8056 2 NOR2X1 $T=1972740 2106160 0 0 $X=1972738 $Y=2105758
X611 4 550 549 8079 2 NOR2X1 $T=1990560 1995280 0 180 $X=1988580 $Y=1989840
X612 4 8215 559 8189 2 NOR2X1 $T=2003760 2146480 0 180 $X=2001780 $Y=2141040
X613 4 8329 570 8332 2 NOR2X1 $T=2032800 2206960 0 0 $X=2032798 $Y=2206558
X614 4 573 8323 8303 2 NOR2X1 $T=2035440 2025520 1 180 $X=2033460 $Y=2025118
X615 4 8352 8373 8393 2 NOR2X1 $T=2044680 2126320 0 0 $X=2044678 $Y=2125918
X616 4 8438 8436 8525 2 NOR2X1 $T=2061840 2136400 0 0 $X=2061838 $Y=2135998
X617 4 8479 8513 8522 2 NOR2X1 $T=2072400 2116240 0 0 $X=2072398 $Y=2115838
X618 4 8522 8525 8540 2 NOR2X1 $T=2075700 2136400 0 0 $X=2075698 $Y=2135998
X619 4 8516 588 8552 2 NOR2X1 $T=2077020 2227120 1 0 $X=2077018 $Y=2221680
X620 4 8566 8591 8587 2 NOR2X1 $T=2089560 2116240 1 0 $X=2089558 $Y=2110800
X621 4 8672 8692 8697 2 NOR2X1 $T=2104740 2126320 1 0 $X=2104738 $Y=2120880
X622 4 8697 8701 8693 2 NOR2X1 $T=2109360 2126320 1 180 $X=2107380 $Y=2125918
X623 4 8671 599 8718 2 NOR2X1 $T=2117940 2217040 1 0 $X=2117938 $Y=2211600
X624 4 8719 8763 8701 2 NOR2X1 $T=2120580 2126320 0 0 $X=2120578 $Y=2125918
X625 4 619 8946 8891 2 NOR2X1 $T=2159520 2015440 1 180 $X=2157540 $Y=2015038
X626 4 8891 8968 8994 2 NOR2X1 $T=2162820 2025520 0 0 $X=2162818 $Y=2025118
X627 4 9014 621 8968 2 NOR2X1 $T=2174040 2015440 0 180 $X=2172060 $Y=2010000
X628 4 8990 9035 9036 2 NOR2X1 $T=2178000 2116240 0 0 $X=2177998 $Y=2115838
X629 4 9057 9036 9017 2 NOR2X1 $T=2182620 2136400 1 180 $X=2180640 $Y=2135998
X630 4 9166 9105 9057 2 NOR2X1 $T=2195820 2136400 1 180 $X=2193840 $Y=2135998
X631 4 9184 9253 9295 2 NOR2X1 $T=2230140 2126320 1 180 $X=2228160 $Y=2125918
X632 4 9280 9360 9331 2 NOR2X1 $T=2249940 2136400 0 0 $X=2249938 $Y=2135998
X633 4 9455 9508 9540 2 NOR2X1 $T=2280300 2146480 0 0 $X=2280298 $Y=2146078
X634 4 9514 9600 9698 2 NOR2X1 $T=2308020 2136400 0 0 $X=2308018 $Y=2135998
X635 4 9540 9698 9687 2 NOR2X1 $T=2309340 2146480 1 0 $X=2309338 $Y=2141040
X636 4 9689 9663 9738 2 NOR2X1 $T=2309340 2166640 0 0 $X=2309338 $Y=2166238
X637 4 9725 661 9806 2 NOR2X1 $T=2333100 1995280 1 0 $X=2333098 $Y=1989840
X638 4 9661 9809 9825 2 NOR2X1 $T=2335080 2126320 0 0 $X=2335078 $Y=2125918
X639 4 9825 9939 10074 2 NOR2X1 $T=2362800 2136400 1 0 $X=2362798 $Y=2130960
X640 4 9873 9861 9939 2 NOR2X1 $T=2366100 2106160 1 180 $X=2364120 $Y=2105758
X641 4 9935 10033 10075 2 NOR2X1 $T=2381280 2116240 0 0 $X=2381278 $Y=2115838
X642 4 10035 10036 10078 2 NOR2X1 $T=2392500 2116240 1 0 $X=2392498 $Y=2110800
X643 4 10078 10075 10142 2 NOR2X1 $T=2393820 2126320 0 0 $X=2393818 $Y=2125918
X644 4 10201 10054 10298 2 NOR2X1 $T=2430780 2116240 0 0 $X=2430778 $Y=2115838
X645 4 10202 10335 10383 2 NOR2X1 $T=2445960 2196880 1 0 $X=2445958 $Y=2191440
X646 4 10435 10314 10461 2 NOR2X1 $T=2463780 2106160 1 0 $X=2463778 $Y=2100720
X647 4 10418 10518 10568 2 NOR2X1 $T=2476320 2096080 0 0 $X=2476318 $Y=2095678
X648 4 10556 10542 10496 2 NOR2X1 $T=2486220 2126320 1 180 $X=2484240 $Y=2125918
X649 4 10568 10461 10609 2 NOR2X1 $T=2497440 2106160 1 0 $X=2497438 $Y=2100720
X650 4 697 10658 700 2 NOR2X1 $T=2506020 1995280 0 0 $X=2506018 $Y=1994878
X651 4 10746 10542 10781 2 NOR2X1 $T=2515920 2116240 0 0 $X=2515918 $Y=2115838
X652 4 10610 10542 10723 2 NOR2X1 $T=2517900 2136400 0 180 $X=2515920 $Y=2130960
X653 4 10298 10683 10782 2 NOR2X1 $T=2521200 2116240 0 0 $X=2521198 $Y=2115838
X654 4 707 708 10792 2 NOR2X1 $T=2523180 2227120 0 0 $X=2523178 $Y=2226718
X655 4 10971 10975 10999 2 NOR2X1 $T=2552220 2055760 0 0 $X=2552218 $Y=2055358
X656 4 10999 10987 10976 2 NOR2X1 $T=2556840 2065840 1 180 $X=2554860 $Y=2065438
X657 4 11043 10542 11059 2 NOR2X1 $T=2568060 2126320 0 0 $X=2568058 $Y=2125918
X658 4 11020 10844 10987 2 NOR2X1 $T=2583240 2055760 1 180 $X=2581260 $Y=2055358
X659 2060 2057 2 4 73 NOR2X2 $T=756360 2217040 0 0 $X=756358 $Y=2216638
X660 2136 2134 2 4 79 NOR2X2 $T=776820 2176720 1 180 $X=773520 $Y=2176318
X661 2133 2196 2 4 782 NOR2X2 $T=790680 2227120 1 180 $X=787380 $Y=2226718
X662 2319 2299 2 4 2353 NOR2X2 $T=825660 2206960 1 0 $X=825658 $Y=2201520
X663 2296 2382 2 4 2397 NOR2X2 $T=828300 2186800 0 0 $X=828298 $Y=2186398
X664 2353 2397 2 4 2384 NOR2X2 $T=831600 2206960 1 180 $X=828300 $Y=2206558
X665 2425 2441 2 4 2422 NOR2X2 $T=841500 2176720 0 180 $X=838200 $Y=2171280
X666 2422 2557 2 4 2537 NOR2X2 $T=859980 2176720 0 180 $X=856680 $Y=2171280
X667 2745 2965 2 4 107 NOR2X2 $T=929280 2186800 1 180 $X=925980 $Y=2186398
X668 107 2892 2 4 113 NOR2X2 $T=938520 2217040 0 0 $X=938518 $Y=2216638
X669 2959 2989 2 4 3057 NOR2X2 $T=947100 2166640 0 0 $X=947098 $Y=2166238
X670 3084 3057 2 4 3117 NOR2X2 $T=957660 2176720 1 0 $X=957658 $Y=2171280
X671 3187 3138 2 4 3145 NOR2X2 $T=976800 2126320 1 0 $X=976798 $Y=2120880
X672 2938 3207 2 4 3226 NOR2X2 $T=988680 2025520 0 180 $X=985380 $Y=2020080
X673 3231 3226 2 4 3199 NOR2X2 $T=988020 2035600 0 0 $X=988018 $Y=2035198
X674 3329 3333 2 4 3231 NOR2X2 $T=1002540 2015440 1 180 $X=999240 $Y=2015038
X675 3562 3553 2 4 3362 NOR2X2 $T=1042140 2196880 0 180 $X=1038840 $Y=2191440
X676 3256 3769 2 4 3737 NOR2X2 $T=1085040 2065840 0 180 $X=1081740 $Y=2060400
X677 4951 5077 2 4 5083 NOR2X2 $T=1349700 2136400 0 0 $X=1349698 $Y=2135998
X678 286 3392 2 4 5230 NOR2X2 $T=1385340 2096080 1 0 $X=1385338 $Y=2090640
X679 479 7255 2 4 7167 NOR2X2 $T=1822920 2015440 0 180 $X=1819620 $Y=2010000
X680 5094 7357 2 4 7324 NOR2X2 $T=1838100 2126320 0 180 $X=1834800 $Y=2120880
X681 7333 7324 2 4 7278 NOR2X2 $T=1836120 2116240 1 0 $X=1836118 $Y=2110800
X682 7356 488 2 4 7323 NOR2X2 $T=1841400 2035600 0 0 $X=1841398 $Y=2035198
X683 7454 7323 2 4 7375 NOR2X2 $T=1854600 2025520 0 0 $X=1854598 $Y=2025118
X684 487 7433 2 4 7351 NOR2X2 $T=1854600 2075920 1 0 $X=1854598 $Y=2070480
X685 5705 7528 2 4 7502 NOR2X2 $T=1869780 2055760 1 180 $X=1866480 $Y=2055358
X686 7587 495 2 4 7563 NOR2X2 $T=1883640 2065840 1 180 $X=1880340 $Y=2065438
X687 7563 7502 2 4 7610 NOR2X2 $T=1884960 2055760 0 0 $X=1884958 $Y=2055358
X688 503 7680 2 4 7588 NOR2X2 $T=1902120 2015440 0 0 $X=1902118 $Y=2015038
X689 7752 7872 2 4 7936 NOR2X2 $T=1943700 2217040 0 0 $X=1943698 $Y=2216638
X690 7895 7865 2 4 7900 NOR2X2 $T=1953600 2116240 1 0 $X=1953598 $Y=2110800
X691 524 527 2 4 7865 NOR2X2 $T=1958220 2106160 0 0 $X=1958218 $Y=2105758
X692 8007 7999 2 4 8023 NOR2X2 $T=1979340 2045680 1 0 $X=1979338 $Y=2040240
X693 594 8608 2 4 8671 NOR2X2 $T=2094180 2206960 0 0 $X=2094178 $Y=2206558
X694 657 9699 2 4 9684 NOR2X2 $T=2310660 2227120 1 180 $X=2307360 $Y=2226718
X695 9750 9684 2 4 9755 NOR2X2 $T=2319900 2227120 1 0 $X=2319898 $Y=2221680
X696 664 9859 2 4 9750 NOR2X2 $T=2341680 2227120 0 180 $X=2338380 $Y=2221680
X697 10227 10232 2 4 10202 NOR2X2 $T=2424180 2196880 0 180 $X=2420880 $Y=2191440
X698 10415 10414 2 4 689 NOR2X2 $T=2460480 2015440 0 0 $X=2460478 $Y=2015038
X699 10444 10462 2 4 10335 NOR2X2 $T=2465760 2196880 1 0 $X=2465758 $Y=2191440
X700 10523 10472 2 4 693 NOR2X2 $T=2483580 2025520 1 0 $X=2483578 $Y=2020080
X701 10724 10682 2 4 697 NOR2X2 $T=2504700 2035600 0 180 $X=2501400 $Y=2030160
X702 10685 10662 2 4 10658 NOR2X2 $T=2505360 2025520 0 180 $X=2502060 $Y=2020080
X703 726 11064 2 4 722 NOR2X2 $T=2570700 2015440 1 180 $X=2567400 $Y=2015038
X704 719 10989 2 4 724 NOR2X2 $T=2570040 1995280 0 0 $X=2570038 $Y=1994878
X705 733 11227 2 4 11154 NOR2X2 $T=2594460 2035600 0 180 $X=2591160 $Y=2030160
X706 730 11092 2 4 11226 NOR2X2 $T=2595120 2025520 1 0 $X=2595118 $Y=2020080
X707 11226 11154 2 4 732 NOR2X2 $T=2598420 1995280 0 0 $X=2598418 $Y=1994878
X708 3937 141 2 4 4298 OR2XL $T=1201200 2186800 0 0 $X=1201198 $Y=2186398
X709 166 164 2 4 253 OR2XL $T=1290300 2227120 1 0 $X=1290298 $Y=2221680
X710 285 276 2 4 5185 OR2XL $T=1373460 2055760 1 0 $X=1373458 $Y=2050320
X711 276 5598 2 4 5615 OR2XL $T=1474440 2035600 0 180 $X=1471800 $Y=2030160
X712 325 337 2 4 5840 OR2XL $T=1512060 2025520 1 0 $X=1512058 $Y=2020080
X713 280 346 2 4 5780 OR2XL $T=1517340 2045680 0 180 $X=1514700 $Y=2040240
X714 311 297 2 4 361 OR2XL $T=1560900 1995280 1 180 $X=1558260 $Y=1994878
X715 375 384 2 4 6302 OR2XL $T=1628880 2206960 1 180 $X=1626240 $Y=2206558
X716 10444 10462 2 4 10432 OR2XL $T=2469720 2176720 1 180 $X=2467080 $Y=2176318
X717 2133 2196 84 2 4 NAND2X2 $T=790680 2217040 1 180 $X=787380 $Y=2216638
X718 2745 2965 108 2 4 NAND2X2 $T=940500 2186800 0 0 $X=940498 $Y=2186398
X719 2804 3088 3058 2 4 NAND2X2 $T=943800 2146480 1 180 $X=940500 $Y=2146078
X720 3063 113 3065 2 4 NAND2X2 $T=954360 2217040 1 180 $X=951060 $Y=2216638
X721 3227 3218 3222 2 4 NAND2X2 $T=986700 2075920 1 0 $X=986698 $Y=2070480
X722 3660 3705 3702 2 4 NAND2X2 $T=1075800 2075920 1 180 $X=1072500 $Y=2075518
X723 270 3381 4913 2 4 NAND2X2 $T=1323300 2146480 0 180 $X=1320000 $Y=2141040
X724 347 378 6285 2 4 NAND2X2 $T=1609740 2196880 1 0 $X=1609738 $Y=2191440
X725 5094 7357 7329 2 4 NAND2X2 $T=1846680 2126320 1 0 $X=1846678 $Y=2120880
X726 488 7356 7328 2 4 NAND2X2 $T=1849320 2035600 0 0 $X=1849318 $Y=2035198
X727 5705 7528 7523 2 4 NAND2X2 $T=1874400 2055760 0 0 $X=1874398 $Y=2055358
X728 503 7680 7566 2 4 NAND2X2 $T=1898820 2025520 1 0 $X=1898818 $Y=2020080
X729 7607 7750 7682 2 4 NAND2X2 $T=1903440 2116240 1 180 $X=1900140 $Y=2115838
X730 508 7746 7690 2 4 NAND2X2 $T=1916640 2106160 0 180 $X=1913340 $Y=2100720
X731 7614 7745 7752 2 4 NAND2X2 $T=1919280 2217040 1 180 $X=1915980 $Y=2216638
X732 7810 7758 7841 2 4 NAND2X2 $T=1934460 2045680 1 0 $X=1934458 $Y=2040240
X733 512 519 7828 2 4 NAND2X2 $T=1935780 2196880 0 0 $X=1935778 $Y=2196478
X734 520 517 7775 2 4 NAND2X2 $T=1945020 2035600 1 0 $X=1945018 $Y=2030160
X735 524 527 7864 2 4 NAND2X2 $T=1951620 2106160 0 180 $X=1948320 $Y=2100720
X736 535 536 7984 2 4 NAND2X2 $T=1966140 2065840 1 0 $X=1966138 $Y=2060400
X737 594 8608 8609 2 4 NAND2X2 $T=2094840 2217040 1 180 $X=2091540 $Y=2216638
X738 9474 9470 9587 2 4 NAND2X2 $T=2269740 2025520 1 0 $X=2269738 $Y=2020080
X739 9699 657 9683 2 4 NAND2X2 $T=2310660 2217040 1 180 $X=2307360 $Y=2216638
X740 10227 10232 10199 2 4 NAND2X2 $T=2424180 2186800 0 180 $X=2420880 $Y=2181360
X741 10415 10414 687 2 4 NAND2X2 $T=2459820 2015440 1 0 $X=2459818 $Y=2010000
X742 730 11092 734 2 4 NAND2X2 $T=2602380 2025520 1 0 $X=2602378 $Y=2020080
X743 2524 4 2537 2451 2 2445 AOI21X4 $T=857340 2206960 1 180 $X=850740 $Y=2206558
X744 5083 4 5085 5023 2 5001 AOI21X4 $T=1356300 2146480 1 180 $X=1349700 $Y=2146078
X745 5460 4 5366 5404 2 5210 AOI21X4 $T=1438140 2075920 0 180 $X=1431540 $Y=2070480
X746 7163 4 7010 7165 2 473 AOI21X4 $T=1797180 2005360 1 0 $X=1797178 $Y=1999920
X747 7278 4 7219 7285 2 7295 AOI21X4 $T=1824900 2116240 1 0 $X=1824898 $Y=2110800
X748 7375 4 7260 7382 2 7431 AOI21X4 $T=1844040 2025520 0 0 $X=1844038 $Y=2025118
X749 7610 4 7591 7631 2 7635 AOI21X4 $T=1892220 2055760 1 0 $X=1892218 $Y=2050320
X750 7900 4 7732 7879 2 7755 AOI21X4 $T=1949640 2116240 0 180 $X=1943040 $Y=2110800
X751 7941 4 7936 7847 2 531 AOI21X4 $T=1953600 2217040 0 0 $X=1953598 $Y=2216638
X752 8994 4 8677 9023 2 9181 AOI21X4 $T=2170740 2025520 0 0 $X=2170738 $Y=2025118
X753 9185 4 9210 9249 2 9251 AOI21X4 $T=2218260 2217040 1 0 $X=2218258 $Y=2211600
X754 9487 4 9755 9771 2 9777 AOI21X4 $T=2321220 2217040 1 0 $X=2321218 $Y=2211600
X755 9806 4 9587 662 2 663 AOI21X4 $T=2333100 1995280 0 0 $X=2333098 $Y=1994878
X756 10015 4 10383 10390 2 10395 AOI21X4 $T=2447940 2186800 0 0 $X=2447938 $Y=2186398
X757 95 4 93 2 2447 AND2X2 $T=829620 2065840 0 0 $X=829618 $Y=2065438
X758 2425 4 2441 2 2514 AND2X2 $T=844140 2176720 1 0 $X=844138 $Y=2171280
X759 2384 4 2537 2 2448 AND2X2 $T=853380 2196880 1 180 $X=850740 $Y=2196478
X760 2617 4 2588 2 2655 AND2X2 $T=875160 2186800 0 0 $X=875158 $Y=2186398
X761 2716 4 2751 2 2739 AND2X2 $T=898920 2136400 0 180 $X=896280 $Y=2130960
X762 2906 4 2928 2 2939 AND2X2 $T=934560 2086000 1 0 $X=934558 $Y=2080560
X763 3110 4 3158 2 3256 AND2X2 $T=969540 2055760 0 0 $X=969538 $Y=2055358
X764 3539 4 3519 2 3483 AND2X2 $T=1040160 2166640 0 180 $X=1037520 $Y=2161200
X765 3681 4 3746 2 3363 AND2X2 $T=1063920 2116240 1 180 $X=1061280 $Y=2115838
X766 3758 4 148 2 3722 AND2X2 $T=1087020 2045680 0 180 $X=1084380 $Y=2040240
X767 148 4 3787 2 3817 AND2X2 $T=1092300 2045680 0 0 $X=1092298 $Y=2045278
X768 348 4 783 2 5889 AND2X2 $T=1527900 2227120 0 0 $X=1527898 $Y=2226718
X769 6302 4 6297 2 6270 AND2X2 $T=1615680 2206960 0 180 $X=1613040 $Y=2201520
X770 6479 4 6517 2 402 AND2X2 $T=1662540 1995280 0 0 $X=1662538 $Y=1994878
X771 6620 4 6714 2 420 AND2X2 $T=1706100 2035600 1 0 $X=1706098 $Y=2030160
X772 7430 4 7374 2 7338 AND2X2 $T=1851300 2005360 1 180 $X=1848660 $Y=2004958
X773 7690 4 7750 2 7744 AND2X2 $T=1916640 2096080 0 0 $X=1916638 $Y=2095678
X774 556 4 553 2 8070 AND2X2 $T=1988580 2227120 1 180 $X=1985940 $Y=2226718
X775 537 4 567 2 8352 AND2X2 $T=2047320 2096080 0 180 $X=2044680 $Y=2090640
X776 8700 4 8512 2 8628 AND2X2 $T=2099460 2025520 0 180 $X=2096820 $Y=2020080
X777 537 4 8670 2 8669 AND2X2 $T=2112660 2075920 1 180 $X=2110020 $Y=2075518
X778 9021 4 8970 2 9044 AND2X2 $T=2183280 2206960 0 180 $X=2180640 $Y=2201520
X779 9282 4 9269 2 9182 AND2X2 $T=2230140 2015440 1 180 $X=2227500 $Y=2015038
X780 9687 4 9494 2 9656 AND2X2 $T=2303400 2146480 0 180 $X=2300760 $Y=2141040
X781 9917 4 9930 2 9914 AND2X2 $T=2355540 2206960 0 180 $X=2352900 $Y=2201520
X782 10074 4 10137 2 10221 AND2X2 $T=2416260 2146480 1 0 $X=2416258 $Y=2141040
X783 3237 2 3222 4 117 NAND2X4 $T=990000 2086000 0 180 $X=985380 $Y=2080560
X784 548 2 543 4 8006 NAND2X4 $T=1983960 2035600 0 180 $X=1979340 $Y=2030160
X785 8116 2 8133 4 555 NAND2X4 $T=1994520 2217040 0 0 $X=1994518 $Y=2216638
X786 2540 2514 2 4 2451 OR2X2 $T=852720 2176720 0 180 $X=850080 $Y=2171280
X787 2590 2610 2 4 2614 OR2X2 $T=872520 2116240 1 0 $X=872518 $Y=2110800
X788 2632 2557 2 4 2617 OR2X2 $T=877800 2176720 1 180 $X=875160 $Y=2176318
X789 2665 2707 2 4 2716 OR2X2 $T=891000 2106160 1 0 $X=890998 $Y=2100720
X790 2789 2801 2 4 2841 OR2X2 $T=906840 2086000 1 0 $X=906838 $Y=2080560
X791 2830 2711 2 4 2843 OR2X2 $T=914760 2055760 0 0 $X=914758 $Y=2055358
X792 71 95 2 4 3064 OR2X2 $T=920040 2025520 0 0 $X=920038 $Y=2025118
X793 3412 3444 2 4 3418 OR2X2 $T=1026960 2156560 0 180 $X=1024320 $Y=2151120
X794 3364 3362 2 4 3414 OR2X2 $T=1032240 2196880 1 180 $X=1029600 $Y=2196478
X795 3541 3486 2 4 3563 OR2X2 $T=1053360 2005360 1 0 $X=1053358 $Y=1999920
X796 152 3815 2 4 3783 OR2X2 $T=1100220 2025520 0 180 $X=1097580 $Y=2020080
X797 195 4599 2 4 4505 OR2X2 $T=1254660 2075920 1 180 $X=1252020 $Y=2075518
X798 93 157 2 4 4696 OR2X2 $T=1275780 2015440 1 0 $X=1275778 $Y=2010000
X799 262 213 2 4 4787 OR2X2 $T=1310760 2126320 1 180 $X=1308120 $Y=2125918
X800 4951 4956 2 4 5107 OR2X2 $T=1330560 2156560 1 0 $X=1330558 $Y=2151120
X801 271 3188 2 4 4994 OR2X2 $T=1331220 2206960 1 0 $X=1331218 $Y=2201520
X802 5040 5076 2 4 4998 OR2X2 $T=1353000 2065840 0 180 $X=1350360 $Y=2060400
X803 5323 3387 2 4 5366 OR2X2 $T=1409100 2075920 1 0 $X=1409098 $Y=2070480
X804 308 255 2 4 5399 OR2X2 $T=1424940 2116240 0 180 $X=1422300 $Y=2110800
X805 308 231 2 4 5396 OR2X2 $T=1424940 2146480 0 180 $X=1422300 $Y=2141040
X806 308 244 2 4 5405 OR2X2 $T=1426260 2166640 1 180 $X=1423620 $Y=2166238
X807 308 213 2 4 5487 OR2X2 $T=1430220 2176720 0 0 $X=1430218 $Y=2176318
X808 308 268 2 4 5554 OR2X2 $T=1432860 2166640 1 0 $X=1432858 $Y=2161200
X809 308 195 2 4 5490 OR2X2 $T=1446720 2106160 0 180 $X=1444080 $Y=2100720
X810 308 289 2 4 5555 OR2X2 $T=1450680 2166640 0 0 $X=1450678 $Y=2166238
X811 308 4469 2 4 5640 OR2X2 $T=1483680 2176720 1 180 $X=1481040 $Y=2176318
X812 308 326 2 4 5819 OR2X2 $T=1502820 2116240 0 0 $X=1502818 $Y=2115838
X813 3667 5889 2 4 5961 OR2X2 $T=1535820 2086000 0 0 $X=1535818 $Y=2085598
X814 4086 6191 2 4 6190 OR2X2 $T=1595880 2045680 0 0 $X=1595878 $Y=2045278
X815 373 381 2 4 6248 OR2X2 $T=1605120 2086000 0 0 $X=1605118 $Y=2085598
X816 373 381 2 4 6256 OR2X2 $T=1615680 2086000 1 180 $X=1613040 $Y=2085598
X817 373 381 2 4 6255 OR2X2 $T=1613700 2106160 1 0 $X=1613698 $Y=2100720
X818 4742 6338 2 4 6329 OR2X2 $T=1623600 2015440 0 0 $X=1623598 $Y=2015038
X819 396 130 2 4 6480 OR2X2 $T=1653300 2035600 0 0 $X=1653298 $Y=2035198
X820 417 6720 2 4 6694 OR2X2 $T=1710060 2005360 1 0 $X=1710058 $Y=1999920
X821 6057 6723 2 4 6721 OR2X2 $T=1710060 2075920 1 0 $X=1710058 $Y=2070480
X822 432 6768 2 4 6764 OR2X2 $T=1719960 2065840 0 180 $X=1717320 $Y=2060400
X823 5362 7030 2 4 6964 OR2X2 $T=1780680 2096080 0 0 $X=1780678 $Y=2095678
X824 465 7080 2 4 7045 OR2X2 $T=1793220 2075920 0 180 $X=1790580 $Y=2070480
X825 7261 5149 2 4 7194 OR2X2 $T=1822260 2106160 0 180 $X=1819620 $Y=2100720
X826 563 561 2 4 8236 OR2X2 $T=2014320 2005360 0 180 $X=2011680 $Y=1999920
X827 8291 565 2 4 8282 OR2X2 $T=2026200 2116240 1 0 $X=2026198 $Y=2110800
X828 578 8405 2 4 8408 OR2X2 $T=2048640 2206960 0 0 $X=2048638 $Y=2206558
X829 8454 581 2 4 8407 OR2X2 $T=2059200 2015440 1 180 $X=2056560 $Y=2015038
X830 8589 587 2 4 8512 OR2X2 $T=2088900 2015440 0 0 $X=2088898 $Y=2015038
X831 602 598 2 4 8700 OR2X2 $T=2110020 2005360 0 180 $X=2107380 $Y=1999920
X832 8829 8808 2 4 8812 OR2X2 $T=2139060 2136400 0 0 $X=2139058 $Y=2135998
X833 8892 8929 2 4 8883 OR2X2 $T=2154240 2136400 0 0 $X=2154238 $Y=2135998
X834 620 8989 2 4 8970 OR2X2 $T=2170080 2206960 1 180 $X=2167440 $Y=2206558
X835 8968 8876 2 4 9066 OR2X2 $T=2172720 2015440 0 0 $X=2172718 $Y=2015038
X836 623 9064 2 4 9021 OR2X2 $T=2183940 2196880 1 0 $X=2183938 $Y=2191440
X837 627 9168 2 4 9210 OR2X2 $T=2204400 2217040 0 0 $X=2204398 $Y=2216638
X838 9215 9295 2 4 9320 OR2X2 $T=2230140 2146480 0 0 $X=2230138 $Y=2146078
X839 637 9273 2 4 9282 OR2X2 $T=2234100 2005360 0 0 $X=2234098 $Y=2004958
X840 9331 9295 2 4 9337 OR2X2 $T=2240700 2146480 1 0 $X=2240698 $Y=2141040
X841 641 9322 2 4 9344 OR2X2 $T=2242020 2217040 1 0 $X=2242018 $Y=2211600
X842 9181 9357 2 4 9474 OR2X2 $T=2246640 2025520 0 0 $X=2246638 $Y=2025118
X843 9245 644 2 4 9356 OR2X2 $T=2254560 2015440 0 0 $X=2254558 $Y=2015038
X844 664 9859 2 4 9830 OR2X2 $T=2345640 2217040 1 0 $X=2345638 $Y=2211600
X845 667 9918 2 4 9917 OR2X2 $T=2356200 2217040 1 180 $X=2353560 $Y=2216638
X846 10225 10290 2 4 10443 OR2X2 $T=2463120 2116240 1 0 $X=2463118 $Y=2110800
X847 10787 10852 2 4 10977 OR2X2 $T=2535060 2075920 0 0 $X=2535058 $Y=2075518
X848 10554 10937 2 4 10943 OR2X2 $T=2546940 2096080 1 0 $X=2546938 $Y=2090640
X849 53 2 4 59 1929 NAND2XL $T=725340 2075920 0 0 $X=725338 $Y=2075518
X850 69 2 4 2076 784 NAND2XL $T=757020 2227120 0 0 $X=757018 $Y=2226718
X851 95 2 4 59 2520 NAND2XL $T=841500 2035600 1 0 $X=841498 $Y=2030160
X852 95 2 4 51 2558 NAND2XL $T=852060 2035600 1 0 $X=852058 $Y=2030160
X853 51 2 4 59 2559 NAND2XL $T=853380 2025520 1 0 $X=853378 $Y=2020080
X854 93 2 4 2885 2983 NAND2XL $T=947100 1995280 1 180 $X=945120 $Y=1994878
X855 3432 2 4 3418 3279 NAND2XL $T=1021680 2166640 0 180 $X=1019700 $Y=2161200
X856 3619 2 4 3482 3437 NAND2XL $T=1050060 2176720 0 180 $X=1048080 $Y=2171280
X857 3861 2 4 3783 3691 NAND2XL $T=1100220 2035600 0 180 $X=1098240 $Y=2030160
X858 4507 2 4 4505 4503 NAND2XL $T=1241460 2075920 1 180 $X=1239480 $Y=2075518
X859 4543 2 4 4535 4531 NAND2XL $T=1246740 2106160 1 180 $X=1244760 $Y=2105758
X860 231 2 4 233 4543 NAND2XL $T=1251360 2106160 0 180 $X=1249380 $Y=2100720
X861 4638 2 4 4541 235 NAND2XL $T=1257300 2227120 0 180 $X=1255320 $Y=2221680
X862 157 2 4 93 4483 NAND2XL $T=1269180 2015440 1 0 $X=1269178 $Y=2010000
X863 4735 2 4 4728 4701 NAND2XL $T=1285680 2116240 0 180 $X=1283700 $Y=2110800
X864 4797 2 4 4787 4695 NAND2XL $T=1294920 2126320 1 180 $X=1292940 $Y=2125918
X865 4728 2 4 4787 4849 NAND2XL $T=1308120 2116240 1 180 $X=1306140 $Y=2115838
X866 213 2 4 262 4797 NAND2XL $T=1310760 2136400 1 180 $X=1308780 $Y=2135998
X867 6257 2 4 6190 6286 NAND2XL $T=1610400 2045680 1 0 $X=1610398 $Y=2040240
X868 384 2 4 375 6297 NAND2XL $T=1620300 2217040 0 180 $X=1618320 $Y=2211600
X869 6335 2 4 6329 6357 NAND2XL $T=1628880 2005360 0 0 $X=1628878 $Y=2004958
X870 130 2 4 396 6481 NAND2XL $T=1653960 2035600 1 0 $X=1653958 $Y=2030160
X871 6697 2 4 6694 6638 NAND2XL $T=1701480 2015440 0 180 $X=1699500 $Y=2010000
X872 6715 2 4 6721 6755 NAND2XL $T=1707420 2065840 0 0 $X=1707418 $Y=2065438
X873 6770 2 4 424 6743 NAND2XL $T=1719960 2045680 0 180 $X=1717980 $Y=2040240
X874 6850 2 4 6764 6823 NAND2XL $T=1743720 2065840 0 180 $X=1741740 $Y=2060400
X875 7047 2 4 7045 7024 NAND2XL $T=1785300 2065840 0 180 $X=1783320 $Y=2060400
X876 7166 2 4 7170 7193 NAND2XL $T=1801800 2116240 0 0 $X=1801798 $Y=2115838
X877 7257 2 4 7194 7173 NAND2XL $T=1822260 2086000 1 180 $X=1820280 $Y=2085598
X878 7592 2 4 7607 7613 NAND2XL $T=1891560 2116240 0 0 $X=1891558 $Y=2115838
X879 7775 2 4 7758 7778 NAND2XL $T=1921920 2035600 1 0 $X=1921918 $Y=2030160
X880 7745 2 4 512 7807 NAND2XL $T=1924560 2196880 0 0 $X=1924558 $Y=2196478
X881 7810 2 4 7788 7782 NAND2XL $T=1926540 2055760 1 180 $X=1924560 $Y=2055358
X882 396 2 4 513 7877 NAND2XL $T=1935120 1995280 0 0 $X=1935118 $Y=1994878
X883 8215 2 4 559 8190 NAND2XL $T=2011680 2146480 0 180 $X=2009700 $Y=2141040
X884 537 2 4 538 8243 NAND2XL $T=2018940 2086000 1 0 $X=2018938 $Y=2080560
X885 568 2 4 566 8290 NAND2XL $T=2029500 2065840 1 0 $X=2029498 $Y=2060400
X886 8439 2 4 8408 8400 NAND2XL $T=2051940 2206960 0 180 $X=2049960 $Y=2201520
X887 8437 2 4 8407 8311 NAND2XL $T=2053260 2045680 0 180 $X=2051280 $Y=2040240
X888 8740 2 4 8700 8607 NAND2XL $T=2125200 2025520 0 180 $X=2123220 $Y=2020080
X889 8823 2 4 8812 8805 NAND2XL $T=2135760 2146480 1 180 $X=2133780 $Y=2146078
X890 8890 2 4 8883 8871 NAND2XL $T=2150280 2166640 0 180 $X=2148300 $Y=2161200
X891 8975 2 4 8970 8927 NAND2XL $T=2164800 2206960 1 180 $X=2162820 $Y=2206558
X892 9037 2 4 9021 8995 NAND2XL $T=2179980 2186800 1 180 $X=2178000 $Y=2186398
X893 9014 2 4 621 8972 NAND2XL $T=2180640 2015440 1 0 $X=2180638 $Y=2010000
X894 9169 2 4 9210 9187 NAND2XL $T=2214300 2217040 1 180 $X=2212320 $Y=2216638
X895 636 2 4 9214 9252 NAND2XL $T=2222880 1995280 1 0 $X=2222878 $Y=1989840
X896 9281 2 4 9257 9246 NAND2XL $T=2226180 2146480 1 180 $X=2224200 $Y=2146078
X897 9342 2 4 9344 9423 NAND2XL $T=2244000 2196880 0 0 $X=2243998 $Y=2196478
X898 9280 2 4 9360 9341 NAND2XL $T=2247300 2136400 1 0 $X=2247298 $Y=2130960
X899 9425 2 4 9356 9302 NAND2XL $T=2255880 2025520 0 180 $X=2253900 $Y=2020080
X900 9455 2 4 9508 9531 NAND2XL $T=2275020 2146480 0 0 $X=2275018 $Y=2146078
X901 9879 2 4 9855 9856 NAND2XL $T=2344980 2146480 0 180 $X=2343000 $Y=2141040
X902 10018 2 4 672 9994 NAND2XL $T=2377980 2217040 1 180 $X=2376000 $Y=2216638
X903 10035 2 4 10036 10139 NAND2XL $T=2397780 2116240 1 0 $X=2397778 $Y=2110800
X904 10136 2 4 10137 10145 NAND2XL $T=2400420 2136400 0 0 $X=2400418 $Y=2135998
X905 10435 2 4 10314 10440 NAND2XL $T=2460480 2106160 1 0 $X=2460478 $Y=2100720
X906 10325 2 4 10443 10419 NAND2XL $T=2465100 2116240 1 180 $X=2463120 $Y=2115838
X907 10322 2 4 10560 10563 NAND2XL $T=2486880 2136400 0 0 $X=2486878 $Y=2135998
X908 10443 2 4 10560 10556 NAND2XL $T=2492160 2126320 1 180 $X=2490180 $Y=2125918
X909 10941 2 4 10943 10849 NAND2XL $T=2543640 2106160 0 180 $X=2541660 $Y=2100720
X910 10980 2 4 10977 11070 NAND2XL $T=2562780 2075920 0 0 $X=2562778 $Y=2075518
X911 10943 2 4 10782 11022 NAND2XL $T=2564760 2116240 0 180 $X=2562780 $Y=2110800
X912 2632 2524 2 4 INVX4 $T=867900 2196880 1 180 $X=865260 $Y=2196478
X913 117 3068 2 4 INVX4 $T=985380 2206960 0 0 $X=985378 $Y=2206558
X914 131 3794 2 4 INVX4 $T=1102860 2005360 0 0 $X=1102858 $Y=2004958
X915 140 152 2 4 INVX4 $T=1131900 1995280 0 180 $X=1129260 $Y=1989840
X916 138 150 2 4 INVX4 $T=1131900 2126320 0 0 $X=1131898 $Y=2125918
X917 5778 218 2 4 INVX4 $T=1495560 2126320 1 180 $X=1492920 $Y=2125918
X918 356 294 2 4 INVX4 $T=1553640 2126320 0 0 $X=1553638 $Y=2125918
X919 5573 375 2 4 INVX4 $T=1594560 2206960 0 180 $X=1591920 $Y=2201520
X920 6164 5656 2 4 INVX4 $T=1601160 2146480 0 180 $X=1598520 $Y=2141040
X921 2679 2614 4 2659 2666 2 AOI21X1 $T=886380 2136400 0 180 $X=883740 $Y=2130960
X922 2841 2888 4 2883 2832 2 AOI21X1 $T=926640 2096080 0 180 $X=924000 $Y=2090640
X923 3064 3062 4 3061 2967 2 AOI21X1 $T=953700 2015440 1 180 $X=951060 $Y=2015038
X924 3186 3227 4 3229 3260 2 AOI21X1 $T=998580 2065840 0 180 $X=995940 $Y=2060400
X925 3449 3431 4 3363 3419 2 AOI21X1 $T=1021680 2116240 1 180 $X=1019040 $Y=2115838
X926 3471 3442 4 3449 3335 2 AOI21X1 $T=1026960 2116240 0 180 $X=1024320 $Y=2110800
X927 3783 3725 4 3780 3720 2 AOI21X1 $T=1093620 2035600 0 180 $X=1090980 $Y=2030160
X928 4720 4730 4 4758 4848 2 AOI21X1 $T=1290300 2106160 1 0 $X=1290298 $Y=2100720
X929 4721 4787 4 4794 4811 2 AOI21X1 $T=1296240 2116240 0 0 $X=1296238 $Y=2115838
X930 4932 4888 4 4906 4865 2 AOI21X1 $T=1318680 2075920 1 180 $X=1316040 $Y=2075518
X931 5015 5081 4 5084 279 2 AOI21X1 $T=1353000 1995280 0 0 $X=1352998 $Y=1994878
X932 276 5509 4 5718 5828 2 AOI21X1 $T=1506120 2196880 1 0 $X=1506118 $Y=2191440
X933 5841 5839 4 5848 5867 2 AOI21X1 $T=1518660 2217040 0 0 $X=1518658 $Y=2216638
X934 6195 6190 4 6189 6056 2 AOI21X1 $T=1597860 2045680 0 180 $X=1595220 $Y=2040240
X935 6334 6329 4 6324 6254 2 AOI21X1 $T=1623600 2005360 0 180 $X=1620960 $Y=1999920
X936 413 6694 4 6709 6710 2 AOI21X1 $T=1707420 2015440 0 180 $X=1704780 $Y=2010000
X937 6761 6721 4 6771 6828 2 AOI21X1 $T=1720620 2075920 1 0 $X=1720618 $Y=2070480
X938 6925 6964 4 6991 7046 2 AOI21X1 $T=1770120 2086000 0 0 $X=1770118 $Y=2085598
X939 7750 7688 4 7686 7589 2 AOI21X1 $T=1904760 2096080 1 180 $X=1902120 $Y=2095678
X940 7758 7772 4 7777 7781 2 AOI21X1 $T=1921260 2045680 1 0 $X=1921258 $Y=2040240
X941 7802 7745 4 7730 7785 2 AOI21X1 $T=1927200 2206960 0 180 $X=1924560 $Y=2201520
X942 8192 8210 4 8209 8208 2 AOI21X1 $T=2008380 2186800 0 180 $X=2005740 $Y=2181360
X943 8236 8206 4 8239 8260 2 AOI21X1 $T=2011020 2025520 1 0 $X=2011018 $Y=2020080
X944 8282 8292 4 8322 8347 2 AOI21X1 $T=2031480 2126320 1 0 $X=2031478 $Y=2120880
X945 8408 8335 4 8473 8519 2 AOI21X1 $T=2061180 2196880 0 0 $X=2061178 $Y=2196478
X946 8540 8404 4 8548 8569 2 AOI21X1 $T=2079000 2136400 0 0 $X=2078998 $Y=2135998
X947 8512 8474 4 8554 8598 2 AOI21X1 $T=2088900 2035600 1 0 $X=2088898 $Y=2030160
X948 589 585 4 8588 8590 2 AOI21X1 $T=2092200 1995280 1 180 $X=2089560 $Y=1994878
X949 8572 8693 4 8694 8717 2 AOI21X1 $T=2104740 2136400 0 0 $X=2104738 $Y=2135998
X950 8554 8700 4 8703 8668 2 AOI21X1 $T=2107380 2015440 0 0 $X=2107378 $Y=2015038
X951 8812 8803 4 8827 8857 2 AOI21X1 $T=2136420 2156560 0 0 $X=2136418 $Y=2156158
X952 8883 8827 4 8930 8926 2 AOI21X1 $T=2155560 2156560 1 0 $X=2155558 $Y=2151120
X953 8987 9021 4 9024 9039 2 AOI21X1 $T=2174040 2206960 1 0 $X=2174038 $Y=2201520
X954 9214 632 4 631 9209 2 AOI21X1 $T=2214300 1995280 1 180 $X=2211660 $Y=1994878
X955 9282 9255 4 9278 9299 2 AOI21X1 $T=2230140 2025520 1 0 $X=2230138 $Y=2020080
X956 9278 9356 4 9453 9470 2 AOI21X1 $T=2264460 2025520 1 0 $X=2264458 $Y=2020080
X957 9494 9230 4 9498 9543 2 AOI21X1 $T=2280960 2156560 1 0 $X=2280958 $Y=2151120
X958 9498 9687 4 9733 9657 2 AOI21X1 $T=2316600 2146480 0 0 $X=2316598 $Y=2146078
X959 10074 9667 4 10140 10143 2 AOI21X1 $T=2400420 2146480 1 0 $X=2400418 $Y=2141040
X960 10140 10142 4 10184 10222 2 AOI21X1 $T=2413620 2126320 0 0 $X=2413618 $Y=2125918
X961 10221 9667 4 10234 10226 2 AOI21X1 $T=2423520 2146480 1 0 $X=2423518 $Y=2141040
X962 9667 10394 4 10412 10416 2 AOI21X1 $T=2453880 2126320 0 0 $X=2453878 $Y=2125918
X963 10486 9667 4 10294 10471 2 AOI21X1 $T=2471040 2136400 0 180 $X=2468400 $Y=2130960
X964 9667 10496 4 10500 10499 2 AOI21X1 $T=2473680 2126320 0 0 $X=2473678 $Y=2125918
X965 10608 10609 4 10655 10684 2 AOI21X1 $T=2499420 2106160 0 0 $X=2499418 $Y=2105758
X966 10657 10590 4 10569 10656 2 AOI21X1 $T=2503380 2136400 0 180 $X=2500740 $Y=2130960
X967 9667 10723 4 10722 10717 2 AOI21X1 $T=2515260 2126320 0 180 $X=2512620 $Y=2120880
X968 10792 701 4 10790 10789 2 AOI21X1 $T=2526480 2217040 1 180 $X=2523840 $Y=2216638
X969 9667 10882 4 10880 714 2 AOI21X1 $T=2541660 2126320 0 180 $X=2539020 $Y=2120880
X970 10886 716 4 10917 10916 2 AOI21X1 $T=2544300 2227120 1 0 $X=2544298 $Y=2221680
X971 10977 11029 4 10973 11094 2 AOI21X1 $T=2575320 2086000 0 0 $X=2575318 $Y=2085598
X972 2790 2717 2 2751 4 2835 OAI21X2 $T=908160 2136400 0 180 $X=902880 $Y=2130960
X973 2976 2967 2 2983 4 2842 OAI21X2 $T=941820 2005360 0 0 $X=941818 $Y=2004958
X974 3166 3068 2 3195 4 3232 OAI21X2 $T=988020 2146480 0 0 $X=988018 $Y=2146078
X975 3362 3433 2 3359 4 3420 OAI21X2 $T=1021680 2196880 0 180 $X=1016400 $Y=2191440
X976 3450 3479 2 3419 4 3388 OAI21X2 $T=1026960 2126320 0 180 $X=1021680 $Y=2120880
X977 3724 3739 2 3720 4 3500 OAI21X2 $T=1082400 2025520 1 180 $X=1077120 $Y=2025118
X978 5019 4951 2 4913 4 5023 OAI21X2 $T=1346400 2146480 1 180 $X=1341120 $Y=2146078
X979 6866 6987 2 6989 4 7021 OAI21X2 $T=1770120 2045680 1 0 $X=1770118 $Y=2040240
X980 7046 7169 2 7187 4 7219 OAI21X2 $T=1801800 2106160 1 0 $X=1801798 $Y=2100720
X981 7296 7323 2 7328 4 7332 OAI21X2 $T=1835460 2025520 1 0 $X=1835458 $Y=2020080
X982 7329 7333 2 7378 4 7285 OAI21X2 $T=1843380 2116240 1 0 $X=1843378 $Y=2110800
X983 7328 7454 2 7374 4 7382 OAI21X2 $T=1850640 2015440 1 180 $X=1845360 $Y=2015038
X984 7523 7563 2 7603 4 7631 OAI21X2 $T=1895520 2065840 0 180 $X=1890240 $Y=2060400
X985 7807 7851 2 7785 4 7812 OAI21X2 $T=1929180 2186800 1 180 $X=1923900 $Y=2186398
X986 519 7752 2 7727 4 7847 OAI21X2 $T=1939740 2217040 1 180 $X=1934460 $Y=2216638
X987 7864 7895 2 7907 4 7879 OAI21X2 $T=1947000 2126320 1 0 $X=1946998 $Y=2120880
X988 7999 7961 2 8006 4 7998 OAI21X2 $T=1966140 2035600 1 0 $X=1966138 $Y=2030160
X989 8006 8007 2 7984 4 8028 OAI21X2 $T=1974060 2045680 0 0 $X=1974058 $Y=2045278
X990 8609 599 2 597 4 604 OAI21X2 $T=2110020 2217040 1 180 $X=2104740 $Y=2216638
X991 9683 9750 2 9796 4 9771 OAI21X2 $T=2327160 2227120 1 0 $X=2327158 $Y=2221680
X992 687 693 2 10522 4 702 OAI21X2 $T=2484900 1995280 0 0 $X=2484898 $Y=1994878
X993 734 11154 2 11250 4 735 OAI21X2 $T=2604360 2005360 1 0 $X=2604358 $Y=1999920
X994 5107 5130 5260 2 4 XNOR2X4 $T=1359600 2156560 1 0 $X=1359598 $Y=2151120
X995 7790 7901 534 2 4 XNOR2X4 $T=1950960 2186800 0 0 $X=1950958 $Y=2186398
X996 9735 9728 655 2 4 XNOR2X4 $T=2319900 2196880 1 180 $X=2308680 $Y=2196478
X997 699 701 10724 2 4 XNOR2X4 $T=2506020 2206960 1 0 $X=2506018 $Y=2201520
X998 3065 2 3068 112 4 111 OAI21X4 $T=956340 2227120 0 180 $X=949080 $Y=2221680
X999 116 2 3068 119 4 785 OAI21X4 $T=976140 2227120 0 0 $X=976138 $Y=2226718
X1000 5004 2 5001 4992 4 273 OAI21X4 $T=1343100 2227120 0 180 $X=1335840 $Y=2221680
X1001 5230 2 5210 5192 4 5085 OAI21X4 $T=1384020 2106160 0 180 $X=1376760 $Y=2100720
X1002 5930 2 5874 5886 4 5460 OAI21X4 $T=1534500 2075920 0 180 $X=1527240 $Y=2070480
X1003 7069 2 7090 7101 4 7010 OAI21X4 $T=1791240 2045680 1 0 $X=1791238 $Y=2040240
X1004 7351 2 7295 7354 4 7260 OAI21X4 $T=1838100 2065840 1 0 $X=1838098 $Y=2060400
X1005 7588 2 7431 7566 4 7591 OAI21X4 $T=1888260 2015440 0 0 $X=1888258 $Y=2015038
X1006 7682 2 7635 7681 4 7732 OAI21X4 $T=1904100 2116240 1 0 $X=1904098 $Y=2110800
X1007 7841 2 7755 7878 4 7962 OAI21X4 $T=1941060 2045680 1 0 $X=1941058 $Y=2040240
X1008 7872 2 7851 519 4 7901 OAI21X4 $T=1950300 2196880 0 180 $X=1943040 $Y=2191440
X1009 9424 2 9251 9457 4 9487 OAI21X4 $T=2259840 2217040 1 0 $X=2259838 $Y=2211600
X1010 9684 2 9655 9683 4 9728 OAI21X4 $T=2311980 2206960 0 0 $X=2311978 $Y=2206558
X1011 9777 2 9996 10011 4 10015 OAI21X4 $T=2372700 2206960 1 0 $X=2372698 $Y=2201520
X1012 333 2 5705 4 CLKBUFX8 $T=1487640 2227120 0 0 $X=1487638 $Y=2226718
X1013 332 2 5321 4 CLKBUFX8 $T=1492920 2106160 1 0 $X=1492918 $Y=2100720
X1014 6389 2 328 4 CLKBUFX8 $T=1638780 2075920 1 180 $X=1634160 $Y=2075518
X1015 6633 2 369 4 CLKBUFX8 $T=1691580 2106160 0 0 $X=1691578 $Y=2105758
X1016 6618 2 414 4 CLKBUFX8 $T=1692240 2065840 1 0 $X=1692238 $Y=2060400
X1017 6746 2 386 4 CLKBUFX8 $T=1723260 2146480 0 0 $X=1723258 $Y=2146078
X1018 6851 2 349 4 CLKBUFX8 $T=1740420 2106160 1 0 $X=1740418 $Y=2100720
X1019 7689 2 504 4 CLKBUFX8 $T=1905420 1995280 0 180 $X=1900800 $Y=1989840
X1020 7729 2 505 4 CLKBUFX8 $T=1913340 2075920 0 180 $X=1908720 $Y=2070480
X1021 7733 2 506 4 CLKBUFX8 $T=1915980 2005360 0 180 $X=1911360 $Y=1999920
X1022 7789 2 511 4 CLKBUFX8 $T=1926540 2075920 0 180 $X=1921920 $Y=2070480
X1023 7938 2 525 4 CLKBUFX8 $T=1955580 2015440 1 180 $X=1950960 $Y=2015038
X1024 617 2 616 4 CLKBUFX8 $T=2159520 2227120 1 180 $X=2154900 $Y=2226718
X1025 2572 2524 4 2 2710 XOR2X2 $T=863280 2206960 1 0 $X=863278 $Y=2201520
X1026 2986 3111 4 2 3140 XOR2X2 $T=958980 2206960 1 0 $X=958978 $Y=2201520
X1027 3206 3068 4 2 3337 XOR2X2 $T=983400 2156560 0 0 $X=983398 $Y=2156158
X1028 3330 3260 4 2 3387 XOR2X2 $T=999240 2075920 1 0 $X=999238 $Y=2070480
X1029 3968 3984 4 2 4108 XOR2X2 $T=1137840 2075920 1 0 $X=1137838 $Y=2070480
X1030 4027 3988 4 2 4086 XOR2X2 $T=1149720 2055760 1 0 $X=1149718 $Y=2050320
X1031 5026 5001 4 2 5094 XOR2X2 $T=1347060 2176720 1 0 $X=1347058 $Y=2171280
X1032 5127 5124 4 2 5149 XOR2X2 $T=1360260 2126320 1 0 $X=1360258 $Y=2120880
X1033 5248 5210 4 2 5362 XOR2X2 $T=1398540 2106160 1 0 $X=1398538 $Y=2100720
X1034 7338 7332 4 2 485 XOR2X2 $T=1840080 1995280 1 180 $X=1833480 $Y=1994878
X1035 7522 7525 4 2 492 XOR2X2 $T=1876380 2035600 0 180 $X=1869780 $Y=2030160
X1036 8995 8992 4 2 618 XOR2X2 $T=2172060 2196880 0 180 $X=2165460 $Y=2191440
X1037 9546 9542 4 2 7455 XOR2X2 $T=2286240 1995280 1 180 $X=2279640 $Y=1994878
X1038 9666 9662 4 2 7680 XOR2X2 $T=2305380 2005360 1 180 $X=2298780 $Y=2004958
X1039 675 674 4 2 7746 XOR2X2 $T=2374680 2005360 0 180 $X=2368080 $Y=1999920
X1040 683 684 4 2 10444 XOR2X2 $T=2434080 2217040 1 0 $X=2434078 $Y=2211600
X1041 151 2 163 4 INVX2 $T=1210440 1995280 1 180 $X=1208460 $Y=1994878
X1042 232 2 234 4 INVX2 $T=1250040 2136400 0 0 $X=1250038 $Y=2135998
X1043 243 2 242 4 INVX2 $T=1270500 2176720 1 0 $X=1270498 $Y=2171280
X1044 256 2 257 4 INVX2 $T=1294260 2156560 1 0 $X=1294258 $Y=2151120
X1045 259 2 260 4 INVX2 $T=1302180 2166640 0 0 $X=1302178 $Y=2166238
X1046 265 2 266 4 INVX2 $T=1312740 2146480 0 0 $X=1312738 $Y=2146078
X1047 276 2 213 4 INVX2 $T=1420320 2227120 0 0 $X=1420318 $Y=2226718
X1048 5783 2 215 4 INVX2 $T=1494900 2096080 1 180 $X=1492920 $Y=2095678
X1049 6018 2 356 4 INVX2 $T=1545720 2146480 0 180 $X=1543740 $Y=2141040
X1050 454 2 476 4 INVX2 $T=1881660 2176720 1 0 $X=1881658 $Y=2171280
X1051 494 2 222 4 INVX2 $T=1882980 2005360 0 0 $X=1882978 $Y=2004958
X1052 7591 2 7525 4 INVX2 $T=1890900 2035600 0 0 $X=1890898 $Y=2035198
X1053 449 2 467 4 INVX2 $T=1896840 2166640 1 0 $X=1896838 $Y=2161200
X1054 451 2 472 4 INVX2 $T=1903440 2186800 0 0 $X=1903438 $Y=2186398
X1055 466 2 475 4 INVX2 $T=1937760 2176720 1 0 $X=1937758 $Y=2171280
X1056 9251 2 9421 4 INVX2 $T=2269740 2196880 0 0 $X=2269738 $Y=2196478
X1057 9777 2 9910 4 INVX2 $T=2349600 2206960 0 180 $X=2347620 $Y=2201520
X1058 73 4 2 2076 INVXL $T=771540 2227120 0 0 $X=771538 $Y=2226718
X1059 4949 4 2 4906 INVXL $T=1329900 2075920 1 180 $X=1328580 $Y=2075518
X1060 4970 4 2 4932 INVXL $T=1336500 2075920 0 0 $X=1336498 $Y=2075518
X1061 213 4 2 5572 INVXL $T=1434180 2156560 1 0 $X=1434178 $Y=2151120
X1062 371 4 2 5509 INVXL $T=1582020 2206960 1 0 $X=1582018 $Y=2201520
X1063 373 4 2 6215 INVXL $T=1584660 2086000 1 0 $X=1584658 $Y=2080560
X1064 328 4 2 6395 INVXL $T=1646700 2106160 1 180 $X=1645380 $Y=2105758
X1065 322 4 2 360 INVXL $T=1700160 2106160 0 0 $X=1700158 $Y=2105758
X1066 309 4 2 428 INVXL $T=1732500 2146480 1 180 $X=1731180 $Y=2146078
X1067 7010 4 2 7040 INVXL $T=1776060 2005360 0 0 $X=1776058 $Y=2004958
X1068 462 4 2 468 INVXL $T=1829520 2217040 1 180 $X=1828200 $Y=2216638
X1069 574 4 2 569 INVXL $T=2036100 1995280 0 180 $X=2034780 $Y=1989840
X1070 8554 4 2 8521 INVXL $T=2080320 2035600 0 180 $X=2079000 $Y=2030160
X1071 8404 4 2 8514 INVXL $T=2080320 2146480 1 180 $X=2079000 $Y=2146078
X1072 625 4 2 9214 INVXL $T=2202420 1995280 1 0 $X=2202418 $Y=1989840
X1073 9295 4 2 9257 INVXL $T=2224200 2146480 0 180 $X=2222880 $Y=2141040
X1074 651 4 2 9603 INVXL $T=2293500 1995280 1 0 $X=2293498 $Y=1989840
X1075 9540 4 2 9654 INVXL $T=2302740 2166640 0 180 $X=2301420 $Y=2161200
X1076 9825 4 2 9855 INVXL $T=2346300 2136400 1 0 $X=2346298 $Y=2130960
X1077 10075 4 2 10137 INVXL $T=2393160 2136400 1 0 $X=2393158 $Y=2130960
X1078 10294 4 2 10320 INVXL $T=2438700 2136400 0 180 $X=2437380 $Y=2130960
X1079 11094 4 2 11140 INVXL $T=2588520 2096080 1 0 $X=2588518 $Y=2090640
X1080 2650 2713 4 2 2745 XNOR2X2 $T=892320 2166640 1 0 $X=892318 $Y=2161200
X1081 2633 2835 4 2 2959 XNOR2X2 $T=915420 2136400 1 0 $X=915418 $Y=2130960
X1082 3114 3139 4 2 3188 XNOR2X2 $T=972180 2196880 1 0 $X=972178 $Y=2191440
X1083 3224 3232 4 2 3381 XNOR2X2 $T=988020 2136400 0 0 $X=988018 $Y=2135998
X1084 3487 3227 4 2 3667 XNOR2X2 $T=1031580 2075920 1 0 $X=1031578 $Y=2070480
X1085 7683 7615 4 2 501 XNOR2X2 $T=1902780 2045680 1 180 $X=1895520 $Y=2045278
X1086 8927 615 4 2 614 XNOR2X2 $T=2155560 2206960 0 180 $X=2148300 $Y=2201520
X1087 8928 8923 4 2 7471 XNOR2X2 $T=2156880 2035600 1 180 $X=2149620 $Y=2035198
X1088 9187 9185 4 2 633 XNOR2X2 $T=2206380 2206960 0 0 $X=2206378 $Y=2206558
X1089 9423 9421 4 2 643 XNOR2X2 $T=2256540 2196880 0 180 $X=2249280 $Y=2191440
X1090 680 681 4 2 7939 XNOR2X2 $T=2409660 2015440 0 180 $X=2402400 $Y=2010000
X1091 93 95 2 4 2358 XOR2X1 $T=819060 2055760 0 0 $X=819058 $Y=2055358
X1092 2719 95 2 4 2741 XOR2X1 $T=893640 2055760 0 0 $X=893638 $Y=2055358
X1093 59 51 2 4 2719 XOR2X1 $T=904200 2025520 0 180 $X=898920 $Y=2020080
X1094 3110 3142 2 4 3255 XOR2X1 $T=966900 2055760 1 0 $X=966898 $Y=2050320
X1095 3278 3271 2 4 2913 XOR2X1 $T=999240 2206960 0 180 $X=993960 $Y=2201520
X1096 3279 3273 2 4 2989 XOR2X1 $T=999900 2166640 0 180 $X=994620 $Y=2161200
X1097 3334 3335 2 4 3088 XOR2X1 $T=1003860 2116240 0 180 $X=998580 $Y=2110800
X1098 3447 3442 2 4 3230 XOR2X1 $T=1025640 2096080 1 180 $X=1020360 $Y=2095678
X1099 3514 3511 2 4 3187 XOR2X1 $T=1038180 2126320 0 180 $X=1032900 $Y=2120880
X1100 3625 3548 2 4 3207 XOR2X1 $T=1056000 2015440 1 180 $X=1050720 $Y=2015038
X1101 3691 3683 2 4 3481 XOR2X1 $T=1071840 2045680 0 180 $X=1066560 $Y=2040240
X1102 3817 3758 2 4 3769 XOR2X1 $T=1100880 2055760 0 180 $X=1095600 $Y=2050320
X1103 3959 3962 2 4 3956 XOR2X1 $T=1137180 2035600 1 180 $X=1131900 $Y=2035198
X1104 3666 125 2 4 4074 XOR2X1 $T=1154340 2186800 0 180 $X=1149060 $Y=2181360
X1105 4531 4534 2 4 230 XOR2X1 $T=1244100 2086000 0 0 $X=1244098 $Y=2085598
X1106 4483 4603 2 4 4637 XOR2X1 $T=1254000 2015440 1 0 $X=1253998 $Y=2010000
X1107 4695 4684 2 4 237 XOR2X1 $T=1278420 2126320 0 180 $X=1273140 $Y=2120880
X1108 252 251 2 4 4599 XOR2X1 $T=1294260 2075920 1 180 $X=1288980 $Y=2075518
X1109 233 4752 2 4 254 XOR2X1 $T=1298880 2005360 1 180 $X=1293600 $Y=2004958
X1110 4866 4865 2 4 261 XOR2X1 $T=1310100 2075920 1 180 $X=1304820 $Y=2075518
X1111 252 262 2 4 267 XOR2X1 $T=1320000 1995280 1 180 $X=1314720 $Y=1994878
X1112 4972 4975 2 4 274 XOR2X1 $T=1333200 2045680 1 0 $X=1333198 $Y=2040240
X1113 5930 5966 2 4 6057 XOR2X1 $T=1547700 2075920 1 0 $X=1547698 $Y=2070480
X1114 6056 6117 2 4 372 XOR2X1 $T=1576080 2045680 0 0 $X=1576078 $Y=2045278
X1115 6866 6946 2 4 6698 XOR2X1 $T=1760880 2035600 1 180 $X=1755600 $Y=2035198
X1116 7041 7040 2 4 6949 XOR2X1 $T=1783320 2015440 1 180 $X=1778040 $Y=2015038
X1117 7074 7069 2 4 6943 XOR2X1 $T=1790580 2045680 1 180 $X=1785300 $Y=2045278
X1118 7193 7209 2 4 7168 XOR2X1 $T=1811700 2086000 0 180 $X=1806420 $Y=2080560
X1119 7301 7295 2 4 484 XOR2X1 $T=1832820 2065840 0 180 $X=1827540 $Y=2060400
X1120 7316 7314 2 4 7189 XOR2X1 $T=1835460 2096080 0 180 $X=1830180 $Y=2090640
X1121 7503 7431 2 4 491 XOR2X1 $T=1869120 2015440 1 180 $X=1863840 $Y=2015038
X1122 7744 7688 2 4 7729 XOR2X1 $T=1916640 2086000 1 180 $X=1911360 $Y=2085598
X1123 7782 7781 2 4 7733 XOR2X1 $T=1925220 2045680 1 180 $X=1919940 $Y=2045278
X1124 521 7873 2 4 522 XOR2X1 $T=1942380 1995280 1 0 $X=1942378 $Y=1989840
X1125 7960 7961 2 4 7938 XOR2X1 $T=1960200 2035600 0 180 $X=1954920 $Y=2030160
X1126 537 538 2 4 8025 XOR2X1 $T=1968780 2075920 0 0 $X=1968778 $Y=2075518
X1127 8001 8055 2 4 545 XOR2X1 $T=1979340 2075920 0 0 $X=1979338 $Y=2075518
X1128 8187 8191 2 4 558 XOR2X1 $T=2005080 2106160 1 180 $X=1999800 $Y=2105758
X1129 8243 8244 2 4 8234 XOR2X1 $T=2015640 2086000 0 180 $X=2010360 $Y=2080560
X1130 8261 8260 2 4 6944 XOR2X1 $T=2018280 2035600 1 180 $X=2013000 $Y=2035198
X1131 567 537 2 4 8291 XOR2X1 $T=2030160 2096080 0 180 $X=2024880 $Y=2090640
X1132 8208 8310 2 4 572 XOR2X1 $T=2030160 2186800 1 0 $X=2030158 $Y=2181360
X1133 8519 8544 2 4 592 XOR2X1 $T=2077680 2196880 0 0 $X=2077678 $Y=2196478
X1134 8607 8598 2 4 7188 XOR2X1 $T=2094180 2035600 1 180 $X=2088900 $Y=2035198
X1135 595 8590 2 4 8589 XOR2X1 $T=2096820 2005360 0 180 $X=2091540 $Y=1999920
X1136 8670 537 2 4 8551 XOR2X1 $T=2102100 2075920 1 180 $X=2096820 $Y=2075518
X1137 8629 8667 2 4 596 XOR2X1 $T=2098140 2196880 1 0 $X=2098138 $Y=2191440
X1138 8676 8673 2 4 8695 XOR2X1 $T=2102100 2166640 0 0 $X=2102098 $Y=2166238
X1139 8788 609 2 4 8946 XOR2X1 $T=2131800 2005360 0 0 $X=2131798 $Y=2004958
X1140 8871 8857 2 4 8851 XOR2X1 $T=2147640 2176720 0 180 $X=2142360 $Y=2171280
X1141 9025 9016 2 4 9011 XOR2X1 $T=2178000 2166640 0 180 $X=2172720 $Y=2161200
X1142 630 9209 2 4 9245 XOR2X1 $T=2209020 2005360 1 0 $X=2209018 $Y=1999920
X1143 9302 9299 2 4 7356 XOR2X1 $T=2235420 2035600 0 180 $X=2230140 $Y=2030160
X1144 9335 9333 2 4 9316 XOR2X1 $T=2243340 2166640 1 180 $X=2238060 $Y=2166238
X1145 9535 9543 2 4 9522 XOR2X1 $T=2284920 2176720 1 180 $X=2279640 $Y=2176318
X1146 9795 9738 2 4 9775 XOR2X1 $T=2332440 2166640 1 180 $X=2327160 $Y=2166238
X1147 10145 10143 2 4 678 XOR2X1 $T=2404380 2156560 1 180 $X=2399100 $Y=2156158
X1148 10220 10226 2 4 10246 XOR2X1 $T=2420880 2156560 1 0 $X=2420878 $Y=2151120
X1149 786 682 2 4 10227 XOR2X1 $T=2432100 2227120 1 180 $X=2426820 $Y=2226718
X1150 10419 10416 2 4 10411 XOR2X1 $T=2460480 2126320 0 180 $X=2455200 $Y=2120880
X1151 10498 10499 2 4 10470 XOR2X1 $T=2476320 2116240 0 180 $X=2471040 $Y=2110800
X1152 10563 10471 2 4 10540 XOR2X1 $T=2489520 2156560 1 180 $X=2484240 $Y=2156158
X1153 10679 10717 2 4 10681 XOR2X1 $T=2512620 2106160 0 180 $X=2507340 $Y=2100720
X1154 710 10789 2 4 712 XOR2X1 $T=2528460 2196880 0 0 $X=2528458 $Y=2196478
X1155 10849 10850 2 4 10815 XOR2X1 $T=2535060 2116240 0 180 $X=2529780 $Y=2110800
X1156 10914 10916 2 4 717 XOR2X1 $T=2544300 2217040 1 0 $X=2544298 $Y=2211600
X1157 11070 11063 2 4 11090 XOR2X1 $T=2575320 2075920 1 0 $X=2575318 $Y=2070480
X1158 2588 4 2557 2572 2 NOR2BX1 $T=867900 2186800 0 180 $X=865260 $Y=2181360
X1159 3494 4 3488 3447 2 NOR2BX1 $T=1034880 2096080 1 180 $X=1032240 $Y=2095678
X1160 125 4 3639 3565 2 NOR2BX1 $T=1056000 2035600 1 0 $X=1055998 $Y=2030160
X1161 3640 4 3565 3625 2 NOR2BX1 $T=1058640 2025520 1 180 $X=1056000 $Y=2025118
X1162 8589 4 8546 8554 2 NOR2BX1 $T=2084280 2015440 1 180 $X=2081640 $Y=2015038
X1163 10443 4 10461 10590 2 NOR2BX1 $T=2494800 2126320 1 0 $X=2494798 $Y=2120880
X1164 10726 4 10658 709 2 NOR2BX1 $T=2525820 1995280 0 0 $X=2525818 $Y=1994878
X1165 10943 4 10972 10974 2 NOR2BX1 $T=2549580 2106160 1 0 $X=2549578 $Y=2100720
X1166 50 52 49 45 4 2 1846 ADDFX2 $T=721380 2045680 0 180 $X=707520 $Y=2040240
X1167 47 51 55 1907 4 2 1999 ADDFX2 $T=710820 2005360 0 0 $X=710818 $Y=2004958
X1168 1870 1871 1887 57 4 2 1910 ADDFX2 $T=711480 2186800 0 0 $X=711478 $Y=2186398
X1169 1869 1872 1888 58 4 2 63 ADDFX2 $T=711480 2227120 1 0 $X=711478 $Y=2221680
X1170 50 49 56 1870 4 2 1945 ADDFX2 $T=713460 2156560 1 0 $X=713458 $Y=2151120
X1171 1951 1956 1945 1930 4 2 1926 ADDFX2 $T=741180 2166640 0 180 $X=727320 $Y=2161200
X1172 59 54 52 1956 4 2 1972 ADDFX2 $T=729300 2116240 1 0 $X=729298 $Y=2110800
X1173 1910 1946 1930 66 4 2 2057 ADDFX2 $T=729960 2206960 0 0 $X=729958 $Y=2206558
X1174 68 65 62 1888 4 2 1946 ADDFX2 $T=745140 2217040 1 180 $X=731280 $Y=2216638
X1175 68 67 64 1887 4 2 1951 ADDFX2 $T=747120 2186800 0 180 $X=733260 $Y=2181360
X1176 52 62 65 2061 4 2 2074 ADDFX2 $T=742500 2136400 1 0 $X=742498 $Y=2130960
X1177 1994 1999 2010 70 4 2 78 ADDFX2 $T=745140 1995280 0 0 $X=745138 $Y=1994878
X1178 1997 2056 1926 2060 4 2 2093 ADDFX2 $T=746460 2186800 0 0 $X=746458 $Y=2186398
X1179 56 72 43 2056 4 2 2058 ADDFX2 $T=764940 2176720 0 180 $X=751080 $Y=2171280
X1180 71 50 53 2098 4 2 2100 ADDFX2 $T=756360 2096080 1 0 $X=756358 $Y=2090640
X1181 2074 2091 2100 2095 4 2 2151 ADDFX2 $T=756360 2116240 0 0 $X=756358 $Y=2115838
X1182 2179 2168 2151 2134 4 2 2133 ADDFX2 $T=786720 2136400 0 180 $X=772860 $Y=2130960
X1183 53 64 68 2168 4 2 2207 ADDFX2 $T=776820 2116240 1 0 $X=776818 $Y=2110800
X1184 49 43 56 2176 4 2 2171 ADDFX2 $T=795960 2176720 0 180 $X=782100 $Y=2171280
X1185 50 71 51 75 4 2 82 ADDFX2 $T=796620 2055760 0 180 $X=782760 $Y=2050320
X1186 47 86 55 2178 4 2 81 ADDFX2 $T=797280 2005360 1 180 $X=783420 $Y=2004958
X1187 55 59 49 2091 4 2 2174 ADDFX2 $T=797280 2075920 1 180 $X=783420 $Y=2075518
X1188 59 54 2209 88 4 2 89 ADDFX2 $T=784080 1995280 0 0 $X=784078 $Y=1994878
X1189 51 71 54 2230 4 2 2224 ADDFX2 $T=787380 2086000 1 0 $X=787378 $Y=2080560
X1190 2171 2210 2224 2211 4 2 2315 ADDFX2 $T=788700 2166640 1 0 $X=788698 $Y=2161200
X1191 95 55 50 2210 4 2 2298 ADDFX2 $T=821700 2075920 0 180 $X=807840 $Y=2070480
X1192 50 68 53 2294 4 2 2424 ADDFX2 $T=809160 2116240 1 0 $X=809158 $Y=2110800
X1193 2362 2352 2298 2318 4 2 2317 ADDFX2 $T=825000 2096080 0 180 $X=811140 $Y=2090640
X1194 65 54 52 2357 4 2 2362 ADDFX2 $T=811800 2106160 0 0 $X=811798 $Y=2105758
X1195 2518 2447 2424 2339 4 2 2402 ADDFX2 $T=848100 2116240 1 180 $X=834240 $Y=2115838
X1196 2358 56 2450 2427 4 2 2571 ADDFX2 $T=836220 2136400 1 0 $X=836218 $Y=2130960
X1197 2421 55 71 2450 4 2 2516 ADDFX2 $T=837540 2055760 0 0 $X=837538 $Y=2055358
X1198 2427 2429 2402 2441 4 2 2560 ADDFX2 $T=839520 2146480 1 0 $X=839518 $Y=2141040
X1199 2421 51 59 2352 4 2 2429 ADDFX2 $T=853380 2086000 0 180 $X=839520 $Y=2080560
X1200 71 59 49 2518 4 2 2522 ADDFX2 $T=840840 2096080 1 0 $X=840838 $Y=2090640
X1201 54 52 2570 2539 4 2 2608 ADDFX2 $T=855360 2106160 0 0 $X=855358 $Y=2105758
X1202 2539 2522 2571 2565 4 2 2630 ADDFX2 $T=855360 2126320 0 0 $X=855358 $Y=2125918
X1203 2516 2631 2608 2603 4 2 2590 ADDFX2 $T=881760 2096080 0 180 $X=867900 $Y=2090640
X1204 55 53 50 2631 4 2 2649 ADDFX2 $T=869220 2055760 1 0 $X=869218 $Y=2050320
X1205 2606 2563 2649 2610 4 2 2665 ADDFX2 $T=871860 2065840 1 0 $X=871858 $Y=2060400
X1206 55 50 2693 2711 4 2 2786 ADDFX2 $T=881760 2005360 0 0 $X=881758 $Y=2004958
X1207 2689 49 2741 2707 4 2 2789 ADDFX2 $T=889020 2075920 1 0 $X=889018 $Y=2070480
X1208 2421 95 71 2689 4 2 2802 ADDFX2 $T=889680 2035600 0 0 $X=889678 $Y=2035198
X1209 2738 54 2802 2801 4 2 2830 ADDFX2 $T=899580 2055760 1 0 $X=899578 $Y=2050320
X1210 3638 3561 3533 3519 4 2 3412 ADDFX2 $T=1050720 2146480 1 180 $X=1036860 $Y=2146078
X1211 3700 133 3663 3553 4 2 3539 ADDFX2 $T=1073160 2156560 0 180 $X=1059300 $Y=2151120
X1212 3766 3694 3661 127 4 2 126 ADDFX2 $T=1075800 2217040 0 180 $X=1061940 $Y=2211600
X1213 131 136 3678 129 4 2 3661 ADDFX2 $T=1076460 2196880 1 180 $X=1062600 $Y=2196478
X1214 140 138 3696 3444 4 2 3681 ADDFX2 $T=1081080 2126320 1 180 $X=1067220 $Y=2125918
X1215 3740 3715 3697 134 4 2 3562 ADDFX2 $T=1081080 2176720 1 180 $X=1067220 $Y=2176318
X1216 3666 141 3748 145 4 2 146 ADDFX2 $T=1076460 2227120 1 0 $X=1076458 $Y=2221680
X1217 139 149 3765 3746 4 2 3626 ADDFX2 $T=1096920 2106160 0 180 $X=1083060 $Y=2100720
X1218 139 132 144 3747 4 2 142 ADDFX2 $T=1096920 2156560 0 180 $X=1083060 $Y=2151120
X1219 3818 151 3747 147 4 2 143 ADDFX2 $T=1102200 2217040 0 180 $X=1088340 $Y=2211600
X1220 157 3818 3794 3698 4 2 3564 ADDFX2 $T=1104840 2096080 0 180 $X=1090980 $Y=2090640
X1221 157 140 3795 3748 4 2 3766 ADDFX2 $T=1104840 2136400 0 180 $X=1090980 $Y=2130960
X1222 157 3815 150 3740 4 2 3663 ADDFX2 $T=1104840 2146480 0 180 $X=1090980 $Y=2141040
X1223 140 3815 159 3847 4 2 154 ADDFX2 $T=1115400 2126320 0 180 $X=1101540 $Y=2120880
X1224 149 164 3847 156 4 2 153 ADDFX2 $T=1115400 2227120 0 180 $X=1101540 $Y=2221680
X1225 3815 131 163 3881 4 2 167 ADDFX2 $T=1104180 2196880 1 0 $X=1104178 $Y=2191440
X1226 4003 3881 3863 160 4 2 155 ADDFX2 $T=1118040 2206960 0 180 $X=1104180 $Y=2201520
X1227 132 125 165 3862 4 2 161 ADDFX2 $T=1120680 2156560 0 180 $X=1106820 $Y=2151120
X1228 138 166 3862 3863 4 2 158 ADDFX2 $T=1120680 2166640 0 180 $X=1106820 $Y=2161200
X1229 125 3937 170 3694 4 2 3697 ADDFX2 $T=1133220 2186800 1 180 $X=1119360 $Y=2186398
X1230 4026 3961 3940 171 4 2 169 ADDFX2 $T=1139160 2227120 0 180 $X=1125300 $Y=2221680
X1231 4006 3696 4077 177 4 2 178 ADDFX2 $T=1145760 2146480 0 0 $X=1145758 $Y=2146078
X1232 180 3561 4074 4026 4 2 4003 ADDFX2 $T=1159620 2186800 1 180 $X=1145760 $Y=2186398
X1233 3666 149 144 4006 4 2 174 ADDFX2 $T=1160940 2136400 1 180 $X=1147080 $Y=2135998
X1234 181 133 4075 176 4 2 3940 ADDFX2 $T=1162920 2217040 1 180 $X=1149060 $Y=2216638
X1235 4125 3638 4156 184 4 2 185 ADDFX2 $T=1169520 2166640 0 0 $X=1169518 $Y=2166238
X1236 3818 141 3561 4140 4 2 4156 ADDFX2 $T=1169520 2176720 0 0 $X=1169518 $Y=2176318
X1237 3937 136 138 4125 4 2 4077 ADDFX2 $T=1184040 2156560 0 180 $X=1170180 $Y=2151120
X1238 4140 150 4167 188 4 2 189 ADDFX2 $T=1172160 2206960 0 0 $X=1172158 $Y=2206558
X1239 138 164 3937 4213 4 2 4205 ADDFX2 $T=1182060 2156560 0 0 $X=1182058 $Y=2156158
X1240 4174 170 4205 198 4 2 199 ADDFX2 $T=1182720 2227120 1 0 $X=1182718 $Y=2221680
X1241 3561 166 136 4323 4 2 4349 ADDFX2 $T=1200540 2156560 1 0 $X=1200538 $Y=2151120
X1242 4296 133 4323 206 4 2 207 ADDFX2 $T=1201200 2206960 0 0 $X=1201198 $Y=2206558
X1243 4213 3795 4349 208 4 2 209 ADDFX2 $T=1203180 2146480 1 0 $X=1203178 $Y=2141040
X1244 163 136 4298 214 4 2 223 ADDFX2 $T=1211760 2196880 1 0 $X=1211758 $Y=2191440
X1245 164 151 181 4541 4 2 4480 ADDFX2 $T=1234860 2217040 1 0 $X=1234858 $Y=2211600
X1246 151 141 180 4486 4 2 225 ADDFX2 $T=1249380 2196880 0 180 $X=1235520 $Y=2191440
X1247 4320 263 262 4851 4 2 4683 ADDFX2 $T=1316700 2106160 0 180 $X=1302840 $Y=2100720
X1248 233 276 4196 5003 4 2 4968 ADDFX2 $T=1353660 2116240 1 180 $X=1339800 $Y=2115838
X1249 215 263 5082 4980 4 2 5040 ADDFX2 $T=1345080 2045680 1 0 $X=1345078 $Y=2040240
X1250 251 280 218 5076 4 2 5074 ADDFX2 $T=1363560 2086000 0 180 $X=1349700 $Y=2080560
X1251 4209 255 5100 5096 4 2 4996 ADDFX2 $T=1367520 2015440 1 180 $X=1353660 $Y=2015038
X1252 244 309 294 5395 4 2 5361 ADDFX2 $T=1432860 2035600 0 180 $X=1419000 $Y=2030160
X1253 310 213 233 313 4 2 5459 ADDFX2 $T=1428240 2055760 1 0 $X=1428238 $Y=2050320
X1254 263 325 322 5597 4 2 318 ADDFX2 $T=1475100 2005360 1 180 $X=1461240 $Y=2004958
X1255 583 8456 538 8436 4 2 8373 ADDFX2 $T=2063160 2106160 1 180 $X=2049300 $Y=2105758
X1256 566 567 584 8479 4 2 8438 ADDFX2 $T=2077680 2096080 0 180 $X=2063820 $Y=2090640
X1257 538 565 8551 8566 4 2 8513 ADDFX2 $T=2072400 2086000 1 0 $X=2072398 $Y=2080560
X1258 584 8456 628 9183 4 2 9165 ADDFX2 $T=2194500 2075920 1 0 $X=2194498 $Y=2070480
X1259 603 647 622 9450 4 2 9513 ADDFX2 $T=2265120 2086000 1 0 $X=2265118 $Y=2080560
X1260 566 649 626 9520 4 2 9456 ADDFX2 $T=2267100 2065840 0 0 $X=2267098 $Y=2065438
X1261 626 622 8704 10138 4 2 10251 ADDFX2 $T=2390520 2086000 0 0 $X=2390518 $Y=2085598
X1262 10756 628 10680 10844 4 2 10852 ADDFX2 $T=2520540 2055760 0 0 $X=2520538 $Y=2055358
X1263 656 647 10881 715 4 2 10975 ADDFX2 $T=2531760 2015440 0 0 $X=2531758 $Y=2015038
X1264 10820 639 10878 10971 4 2 11020 ADDFX2 $T=2539680 2055760 1 0 $X=2539678 $Y=2050320
X1265 2441 2425 2 4 2616 XNOR2X1 $T=844140 2176720 0 0 $X=844138 $Y=2176318
X1266 2603 2630 2 4 2650 XNOR2X1 $T=875160 2156560 0 0 $X=875158 $Y=2156158
X1267 2739 2717 2 4 2804 XNOR2X1 $T=896940 2146480 1 0 $X=896938 $Y=2141040
X1268 2935 2939 2 4 3138 XNOR2X1 $T=934560 2106160 0 0 $X=934558 $Y=2105758
X1269 2945 2834 2 4 2977 XNOR2X1 $T=937860 2086000 0 0 $X=937858 $Y=2085598
X1270 3106 3062 2 4 3122 XNOR2X1 $T=958980 2035600 1 0 $X=958978 $Y=2030160
X1271 3437 3436 2 4 2965 XNOR2X1 $T=1023000 2176720 1 180 $X=1017720 $Y=2176318
X1272 3462 3466 2 4 3333 XNOR2X1 $T=1028280 2005360 1 180 $X=1023000 $Y=2004958
X1273 3509 3500 2 4 3416 XNOR2X1 $T=1037520 2015440 1 180 $X=1032240 $Y=2015038
X1274 141 3937 2 4 4296 XNOR2X1 $T=1199880 2196880 1 0 $X=1199878 $Y=2191440
X1275 139 3987 2 4 4321 XNOR2X1 $T=1203180 2015440 0 0 $X=1203178 $Y=2015038
X1276 4503 4504 2 4 224 XNOR2X1 $T=1241460 2086000 1 180 $X=1236180 $Y=2085598
X1277 4701 4702 2 4 238 XNOR2X1 $T=1280400 2116240 0 180 $X=1275120 $Y=2110800
X1278 4890 4888 2 4 250 XNOR2X1 $T=1314720 2075920 0 180 $X=1309440 $Y=2070480
X1279 276 285 2 4 5100 XNOR2X1 $T=1377420 2035600 1 180 $X=1372140 $Y=2035198
X1280 787 299 2 4 5323 XNOR2X1 $T=1398540 2227120 0 0 $X=1398538 $Y=2226718
X1281 5598 276 2 4 5616 XNOR2X1 $T=1463880 2035600 1 0 $X=1463878 $Y=2030160
X1282 5460 5437 2 4 5741 XNOR2X1 $T=1469160 2075920 1 0 $X=1469158 $Y=2070480
X1283 337 325 2 4 5690 XNOR2X1 $T=1500840 2035600 1 180 $X=1495560 $Y=2035198
X1284 346 280 2 4 5638 XNOR2X1 $T=1519980 2055760 0 180 $X=1514700 $Y=2050320
X1285 297 311 2 4 359 XNOR2X1 $T=1544400 1995280 0 0 $X=1544398 $Y=1994878
X1286 5977 6051 2 4 6080 XNOR2X1 $T=1560900 2086000 1 0 $X=1560898 $Y=2080560
X1287 380 379 2 4 6191 XNOR2X1 $T=1606440 2227120 0 180 $X=1601160 $Y=2221680
X1288 6195 6286 2 4 390 XNOR2X1 $T=1610400 2025520 1 0 $X=1610398 $Y=2020080
X1289 6334 6357 2 4 387 XNOR2X1 $T=1628880 2005360 1 0 $X=1628878 $Y=1999920
X1290 7024 7021 2 4 6931 XNOR2X1 $T=1780020 2055760 1 180 $X=1774740 $Y=2055358
X1291 459 460 2 4 6947 XNOR2X1 $T=1785960 1995280 0 180 $X=1780680 $Y=1989840
X1292 7058 7056 2 4 6948 XNOR2X1 $T=1788600 2005360 0 180 $X=1783320 $Y=1999920
X1293 7091 7173 2 4 7080 XNOR2X1 $T=1806420 2086000 1 180 $X=1801140 $Y=2085598
X1294 7368 7365 2 4 7255 XNOR2X1 $T=1847340 2096080 0 180 $X=1842060 $Y=2090640
X1295 7778 7772 2 4 7689 XNOR2X1 $T=1924560 2025520 0 180 $X=1919280 $Y=2020080
X1296 7830 7829 2 4 7789 XNOR2X1 $T=1937100 2106160 1 180 $X=1931820 $Y=2105758
X1297 7982 7998 2 4 532 XNOR2X1 $T=1968780 2025520 0 180 $X=1963500 $Y=2020080
X1298 8206 8194 2 4 6723 XNOR2X1 $T=2006400 2055760 1 180 $X=2001120 $Y=2055358
X1299 8192 8235 2 4 562 XNOR2X1 $T=2009040 2166640 1 0 $X=2009038 $Y=2161200
X1300 8292 8288 2 4 8278 XNOR2X1 $T=2026200 2126320 1 180 $X=2020920 $Y=2125918
X1301 8311 8307 2 4 7030 XNOR2X1 $T=2031480 2055760 1 180 $X=2026200 $Y=2055358
X1302 8337 571 2 4 8323 XNOR2X1 $T=2036760 2005360 1 180 $X=2031480 $Y=2004958
X1303 8335 8400 2 4 580 XNOR2X1 $T=2047320 2196880 1 0 $X=2047318 $Y=2191440
X1304 8495 8474 2 4 7261 XNOR2X1 $T=2069100 2035600 1 180 $X=2063820 $Y=2035198
X1305 8510 585 2 4 8454 XNOR2X1 $T=2073060 1995280 1 180 $X=2067780 $Y=1994878
X1306 8478 8511 2 4 8515 XNOR2X1 $T=2071740 2156560 1 0 $X=2071738 $Y=2151120
X1307 8741 8720 2 4 600 XNOR2X1 $T=2117940 2206960 0 180 $X=2112660 $Y=2201520
X1308 8747 8745 2 4 605 XNOR2X1 $T=2117940 2156560 0 0 $X=2117938 $Y=2156158
X1309 8805 8803 2 4 8784 XNOR2X1 $T=2133780 2156560 1 180 $X=2128500 $Y=2156158
X1310 8824 8677 2 4 7357 XNOR2X1 $T=2137740 2035600 0 180 $X=2132460 $Y=2030160
X1311 612 8849 2 4 9014 XNOR2X1 $T=2143020 1995280 0 0 $X=2143018 $Y=1994878
X1312 9085 9082 2 4 9108 XNOR2X1 $T=2191200 2156560 0 0 $X=2191198 $Y=2156158
X1313 9182 9181 2 4 7433 XNOR2X1 $T=2207040 2035600 1 180 $X=2201760 $Y=2035198
X1314 9246 9230 2 4 9190 XNOR2X1 $T=2222220 2166640 0 180 $X=2216940 $Y=2161200
X1315 9252 632 2 4 9273 XNOR2X1 $T=2223540 2005360 1 0 $X=2223538 $Y=1999920
X1316 660 9783 2 4 9454 XNOR2X1 $T=2332440 2015440 0 180 $X=2327160 $Y=2010000
X1317 9856 9667 2 4 9878 XNOR2X1 $T=2343000 2156560 1 0 $X=2342998 $Y=2151120
X1318 9929 9928 2 4 9916 XNOR2X1 $T=2358840 2146480 1 180 $X=2353560 $Y=2146078
X1319 669 668 2 4 9909 XNOR2X1 $T=2360820 1995280 1 180 $X=2355540 $Y=1994878
X1320 210 332 2 308 4 218 5711 5689 OAI221XL $T=1488300 2106160 1 0 $X=1488298 $Y=2100720
X1321 217 332 2 308 4 215 5719 5693 OAI221XL $T=1491600 2065840 1 0 $X=1491598 $Y=2060400
X1322 5894 5934 2 251 4 5656 5954 5858 OAI221XL $T=1539780 2166640 1 0 $X=1539778 $Y=2161200
X1323 194 5808 2 308 4 4196 5941 5950 OAI221XL $T=1547040 2116240 1 180 $X=1542420 $Y=2115838
X1324 351 353 2 353 4 6012 5980 358 OAI221XL $T=1554960 2227120 0 180 $X=1550340 $Y=2221680
X1325 197 5808 2 308 4 370 6478 6358 OAI221XL $T=1650000 2146480 0 0 $X=1649998 $Y=2146078
X1326 421 5808 2 308 4 422 6757 6713 OAI221XL $T=1712700 2186800 0 0 $X=1712698 $Y=2186398
X1327 426 5808 2 308 4 293 6791 6724 OAI221XL $T=1720620 2186800 0 0 $X=1720618 $Y=2186398
X1328 429 5808 2 308 4 322 6834 6712 OAI221XL $T=1733820 2166640 1 0 $X=1733818 $Y=2161200
X1329 221 5808 2 308 4 227 6835 6695 OAI221XL $T=1733820 2176720 0 0 $X=1733818 $Y=2176318
X1330 431 5808 2 308 4 310 6857 6867 OAI221XL $T=1739100 2186800 0 0 $X=1739098 $Y=2186398
X1331 436 5808 2 308 4 309 6882 6864 OAI221XL $T=1744380 2156560 0 0 $X=1744378 $Y=2156158
X1332 439 5808 2 308 4 430 6897 6860 OAI221XL $T=1746360 2186800 0 0 $X=1746358 $Y=2186398
X1333 49 1872 52 4 2 42 ADDHXL $T=721380 2217040 0 180 $X=714120 $Y=2211600
X1334 53 788 56 4 2 789 ADDHXL $T=717420 2227120 0 0 $X=717418 $Y=2226718
X1335 54 1871 53 4 2 1869 ADDHXL $T=724680 2176720 1 180 $X=717420 $Y=2176318
X1336 93 2297 47 4 2 2209 ADDHXL $T=823680 2005360 0 180 $X=816420 $Y=1999920
X1337 93 2563 51 4 2 2570 ADDHXL $T=857340 2075920 1 0 $X=857338 $Y=2070480
X1338 93 2693 2421 4 2 2738 ADDHXL $T=890340 1995280 0 0 $X=890338 $Y=1994878
X1339 51 2885 59 4 2 2828 ADDHXL $T=928620 2005360 0 180 $X=921360 $Y=1999920
X1340 130 3533 132 4 2 3700 ADDHXL $T=1062600 2146480 0 0 $X=1062598 $Y=2146078
X1341 130 3639 3666 4 2 3569 ADDHXL $T=1071180 2065840 0 180 $X=1063920 $Y=2060400
X1342 130 3715 139 4 2 3678 ADDHXL $T=1071840 2176720 1 0 $X=1071838 $Y=2171280
X1343 252 5229 285 4 2 5383 ADDHXL $T=1387320 2015440 1 0 $X=1387318 $Y=2010000
X1344 608 8804 537 4 2 8852 ADDHXL $T=2128500 2086000 0 0 $X=2128498 $Y=2085598
X1345 603 9821 647 4 2 9912 ADDHXL $T=2332440 2045680 0 0 $X=2332438 $Y=2045278
X1346 603 9976 649 4 2 10013 ADDHXL $T=2389860 2045680 0 180 $X=2382600 $Y=2040240
X1347 608 10046 647 4 2 10160 ADDHXL $T=2412960 2055760 0 180 $X=2405700 $Y=2050320
X1348 634 10393 649 4 2 10473 ADDHXL $T=2455200 2065840 1 0 $X=2455198 $Y=2060400
X1349 639 10274 656 4 2 10410 ADDHXL $T=2475000 2086000 0 0 $X=2474998 $Y=2085598
X1350 649 10756 647 4 2 10820 ADDHXL $T=2523180 2055760 1 0 $X=2523178 $Y=2050320
X1351 656 10878 649 4 2 10881 ADDHXL $T=2535060 2025520 1 0 $X=2535058 $Y=2020080
X1352 4 93 51 3144 2 NOR2XL $T=963600 2065840 1 0 $X=963598 $Y=2060400
X1353 4 233 4752 4734 2 NOR2XL $T=1290960 2005360 1 180 $X=1288980 $Y=2004958
X1354 4 233 251 4765 2 NOR2XL $T=1290300 2045680 0 0 $X=1290298 $Y=2045278
X1355 4 396 513 7869 2 NOR2XL $T=1925880 1995280 1 0 $X=1925878 $Y=1989840
X1356 4 568 566 8306 2 NOR2XL $T=2030160 2075920 0 180 $X=2028180 $Y=2070480
X1357 4 10298 10230 10394 2 NOR2XL $T=2453220 2136400 0 0 $X=2453218 $Y=2135998
X1358 4 10982 10542 10882 2 NOR2XL $T=2554200 2126320 1 180 $X=2552220 $Y=2125918
X1359 4 11022 10542 11066 2 NOR2XL $T=2565420 2116240 0 0 $X=2565418 $Y=2115838
X1360 4 10987 11065 11091 2 NOR2XL $T=2575320 2096080 1 0 $X=2575318 $Y=2090640
X1361 4 11133 10542 11165 2 NOR2XL $T=2589180 2126320 0 0 $X=2589178 $Y=2125918
X1362 1999 1994 2010 2 4 76 XOR3X2 $T=747120 2015440 1 0 $X=747118 $Y=2010000
X1363 53 54 59 2 4 2015 XOR3X2 $T=760980 2075920 1 180 $X=749100 $Y=2075518
X1364 2842 2786 2828 2 4 2938 XOR3X2 $T=924660 2005360 0 0 $X=924658 $Y=2004958
X1365 4660 4683 4703 2 4 249 XOR3X2 $T=1269840 2086000 1 0 $X=1269838 $Y=2080560
X1366 5015 4996 4980 2 4 272 XOR3X2 $T=1347060 2005360 1 180 $X=1335180 $Y=2004958
X1367 8404 8436 8438 2 4 8398 XOR3X2 $T=2064480 2146480 1 180 $X=2052600 $Y=2146078
X1368 4728 4702 4 4721 2 4684 AOI21XL $T=1283700 2116240 1 180 $X=1281060 $Y=2115838
X1369 4954 4888 4 4965 2 4975 AOI21XL $T=1330560 2075920 1 0 $X=1330558 $Y=2070480
X1370 7194 7091 4 7211 2 7209 AOI21XL $T=1809060 2086000 0 0 $X=1809058 $Y=2085598
X1371 10443 10657 4 10608 2 10562 AOI21XL $T=2503380 2126320 0 180 $X=2500740 $Y=2120880
X1372 9667 10781 4 10847 2 10850 AOI21XL $T=2531100 2116240 0 0 $X=2531098 $Y=2115838
X1373 10973 10976 4 10978 2 10981 AOI21XL $T=2552220 2075920 1 0 $X=2552218 $Y=2070480
X1374 10974 10727 4 10984 2 10990 AOI21XL $T=2553540 2106160 0 0 $X=2553538 $Y=2105758
X1375 10943 10727 4 11029 2 11026 AOI21XL $T=2564760 2106160 0 0 $X=2564758 $Y=2105758
X1376 9667 11059 4 11060 2 11062 AOI21XL $T=2572020 2126320 1 0 $X=2572018 $Y=2120880
X1377 9667 11066 4 11001 2 11063 AOI21XL $T=2577960 2116240 1 180 $X=2575320 $Y=2115838
X1378 11091 10727 4 11110 2 11095 AOI21XL $T=2583240 2106160 0 180 $X=2580600 $Y=2100720
X1379 11155 10727 4 11140 2 11129 AOI21XL $T=2593800 2106160 0 180 $X=2591160 $Y=2100720
X1380 9667 11165 4 11160 2 11175 AOI21XL $T=2596440 2116240 0 0 $X=2596438 $Y=2115838
X1381 3418 3388 3432 2 3436 4 OAI2BB1X1 $T=1019040 2176720 1 0 $X=1019038 $Y=2171280
X1382 351 353 5920 2 5848 4 OAI2BB1X1 $T=1537800 2217040 0 0 $X=1537798 $Y=2216638
X1383 8925 8677 8876 2 8923 4 OAI2BB1X1 $T=2154240 2035600 0 180 $X=2150940 $Y=2030160
X1384 9338 9404 9341 2 9498 4 OAI2BB1X1 $T=2249280 2146480 0 0 $X=2249278 $Y=2146078
X1385 9734 9587 659 2 9783 4 OAI2BB1X1 $T=2319900 2005360 1 0 $X=2319898 $Y=1999920
X1386 9667 9855 9879 2 9928 4 OAI2BB1X1 $T=2348940 2146480 1 0 $X=2348938 $Y=2141040
X1387 10137 10140 10136 2 10234 4 OAI2BB1X1 $T=2407680 2136400 0 0 $X=2407678 $Y=2135998
X1388 10015 10276 10199 2 10317 4 OAI2BB1X1 $T=2440020 2186800 0 0 $X=2440018 $Y=2186398
X1389 2353 2 2337 4 92 NAND2BXL $T=817740 2206960 1 180 $X=815100 $Y=2206558
X1390 3443 2 3366 4 3334 NAND2BXL $T=1010460 2116240 0 180 $X=1007820 $Y=2110800
X1391 3486 2 3461 4 3462 NAND2BXL $T=1026960 2005360 0 180 $X=1024320 $Y=1999920
X1392 4382 2 4443 4 4603 NAND2BXL $T=1242780 2015440 0 0 $X=1242778 $Y=2015038
X1393 5078 2 5126 4 278 NAND2BXL $T=1362240 1995280 0 180 $X=1359600 $Y=1989840
X1394 304 2 335 4 5800 NAND2BXL $T=1505460 2217040 1 0 $X=1505458 $Y=2211600
X1395 378 2 334 4 5426 NAND2BXL $T=1560900 2176720 1 180 $X=1558260 $Y=2176318
X1396 368 2 363 4 6079 NAND2BXL $T=1574100 2196880 1 180 $X=1571460 $Y=2196478
X1397 6099 2 233 4 6052 NAND2BXL $T=1575420 2166640 0 180 $X=1572780 $Y=2161200
X1398 6763 2 6743 4 6717 NAND2BXL $T=1714020 2045680 0 180 $X=1711380 $Y=2040240
X1399 6987 2 6989 4 6946 NAND2BXL $T=1772760 2035600 1 180 $X=1770120 $Y=2035198
X1400 7068 2 7059 4 7041 NAND2BXL $T=1789260 2015440 1 180 $X=1786620 $Y=2015038
X1401 7090 2 7101 4 7074 NAND2BXL $T=1806420 2045680 0 0 $X=1806418 $Y=2045278
X1402 7333 2 7378 4 7368 NAND2BXL $T=1851960 2106160 0 180 $X=1849320 $Y=2100720
X1403 7502 2 7523 4 7522 NAND2BXL $T=1874400 2045680 1 180 $X=1871760 $Y=2045278
X1404 7999 2 8006 4 7960 NAND2BXL $T=1976700 2035600 0 180 $X=1974060 $Y=2030160
X1405 8056 2 8057 4 8055 NAND2BXL $T=1980660 2106160 1 0 $X=1980658 $Y=2100720
X1406 8079 2 547 4 8021 NAND2BXL $T=1987920 1995280 1 180 $X=1985280 $Y=1994878
X1407 8522 2 8493 4 8478 NAND2BXL $T=2068440 2126320 1 180 $X=2065800 $Y=2125918
X1408 8587 2 8584 4 8571 NAND2BXL $T=2088900 2136400 0 180 $X=2086260 $Y=2130960
X1409 599 2 597 4 8741 NAND2BXL $T=2117940 2217040 0 0 $X=2117938 $Y=2216638
X1410 610 2 606 4 8788 NAND2BXL $T=2131140 1995280 1 180 $X=2128500 $Y=1994878
X1411 9036 2 9018 4 9016 NAND2BXL $T=2175360 2156560 1 180 $X=2172720 $Y=2156158
X1412 9057 2 9098 4 9085 NAND2BXL $T=2195160 2146480 1 180 $X=2192520 $Y=2146078
X1413 9331 2 9341 4 9335 NAND2BXL $T=2245320 2156560 1 180 $X=2242680 $Y=2156158
X1414 9540 2 9531 4 9535 NAND2BXL $T=2283600 2166640 0 180 $X=2280960 $Y=2161200
X1415 9698 2 9700 4 9795 NAND2BXL $T=2329800 2146480 0 0 $X=2329798 $Y=2146078
X1416 9939 2 9938 4 9929 NAND2BXL $T=2362140 2116240 1 180 $X=2359500 $Y=2115838
X1417 10568 2 10570 4 10679 NAND2BXL $T=2502060 2106160 1 0 $X=2502058 $Y=2100720
X1418 6143 5719 2 4 CLKBUFX3 $T=1583340 2065840 0 0 $X=1583338 $Y=2065438
X1419 399 6440 2 4 CLKBUFX3 $T=1695540 1995280 1 0 $X=1695538 $Y=1989840
X1420 530 7941 2 4 CLKBUFX3 $T=1954260 2217040 1 0 $X=1954258 $Y=2211600
X1421 240 5321 259 301 4 2 5345 AOI2BB2X1 $T=1399200 2166640 0 0 $X=1399198 $Y=2166238
X1422 216 5321 243 301 4 2 5339 AOI2BB2X1 $T=1401180 2176720 0 0 $X=1401178 $Y=2176318
X1423 205 5321 232 301 4 2 5358 AOI2BB2X1 $T=1406460 2146480 1 0 $X=1406458 $Y=2141040
X1424 258 5321 281 301 4 2 5442 AOI2BB2X1 $T=1409760 2106160 0 0 $X=1409758 $Y=2105758
X1425 200 5321 291 301 4 2 5492 AOI2BB2X1 $T=1410420 2086000 0 0 $X=1410418 $Y=2085598
X1426 202 5808 342 301 4 2 5823 AOI2BB2X1 $T=1510080 2106160 0 0 $X=1510078 $Y=2105758
X1427 1908 1928 1845 60 4 2 61 ADDFHX1 $T=721380 2025520 0 0 $X=721378 $Y=2025118
X1428 2098 2058 1972 1997 4 2 2055 ADDFHX1 $T=765600 2156560 1 180 $X=750420 $Y=2156158
X1429 2061 2095 2055 2097 4 2 2136 ADDFHX1 $T=755040 2146480 1 0 $X=755038 $Y=2141040
X1430 2230 2207 2174 2179 4 2 2175 ADDFHX1 $T=799260 2096080 0 180 $X=784080 $Y=2090640
X1431 2176 2211 2175 2196 4 2 2319 ADDFHX1 $T=785400 2196880 1 0 $X=785398 $Y=2191440
X1432 1886 2 1929 4 1924 1908 NAND3X1 $T=727980 2065840 0 0 $X=727978 $Y=2065438
X1433 2520 2 2558 4 2559 2606 NAND3X1 $T=858660 2035600 1 0 $X=858658 $Y=2030160
X1434 5358 2 5397 4 5396 5400 NAND3X1 $T=1420980 2146480 0 0 $X=1420978 $Y=2146078
X1435 5426 2 5345 4 5405 5406 NAND3X1 $T=1426260 2176720 1 180 $X=1423620 $Y=2176318
X1436 149 151 133 4174 2 4 4167 CMPR32X1 $T=1172820 2217040 1 0 $X=1172818 $Y=2211600
X1437 584 8456 622 8997 2 4 8881 CMPR32X1 $T=2183940 2096080 0 180 $X=2170080 $Y=2090640
X1438 565 608 639 9521 2 4 9599 CMPR32X1 $T=2267100 2075920 1 0 $X=2267098 $Y=2070480
X1439 608 647 626 10392 2 4 10391 CMPR32X1 $T=2442000 2055760 0 0 $X=2441998 $Y=2055358
X1440 3250 3254 3392 3254 3250 2 4 OAI2BB2X2 $T=993300 2045680 0 0 $X=993298 $Y=2045278
X1441 3432 3469 3433 2 3483 4 AOI2BB1X2 $T=1027620 2176720 0 0 $X=1027618 $Y=2176318
X1442 3935 3959 3918 2 3919 4 AOI2BB1X2 $T=1128600 2035600 0 180 $X=1123980 $Y=2030160
X1443 1907 1846 46 44 4 2 1845 ADDFHX2 $T=729960 2015440 1 180 $X=707520 $Y=2015038
X1444 75 2073 2015 1928 4 2 2010 ADDFHX2 $T=770220 2035600 1 180 $X=747780 $Y=2035198
X1445 49 87 2178 1994 4 2 83 ADDFHX2 $T=806520 2015440 0 180 $X=784080 $Y=2010000
X1446 2294 2339 2317 2382 4 2 2425 ADDFHX2 $T=805860 2146480 1 0 $X=805858 $Y=2141040
X1447 2297 2073 82 96 4 2 98 ADDFHX2 $T=807840 2025520 0 0 $X=807838 $Y=2025118
X1448 2357 2318 2315 2299 4 2 2296 ADDFHX2 $T=830280 2176720 0 180 $X=807840 $Y=2171280
X1449 564 8263 2 4 8210 OR2X1 $T=2020920 2176720 0 0 $X=2020918 $Y=2176318
X1450 9057 9018 2 4 9043 OR2X1 $T=2183280 2146480 0 180 $X=2180640 $Y=2141040
X1451 2831 4 2717 2 CLKINVX3 $T=914100 2146480 1 180 $X=912120 $Y=2146078
X1452 115 4 119 2 CLKINVX3 $T=969540 2227120 0 0 $X=969538 $Y=2226718
X1453 3388 4 3273 2 CLKINVX3 $T=1005840 2176720 0 180 $X=1003860 $Y=2171280
X1454 3532 4 3227 2 CLKINVX3 $T=1037520 2065840 0 180 $X=1035540 $Y=2060400
X1455 3918 4 3758 2 CLKINVX3 $T=1110780 2035600 1 180 $X=1108800 $Y=2035198
X1456 3795 4 133 2 CLKINVX3 $T=1135200 2136400 0 0 $X=1135198 $Y=2135998
X1457 157 4 3958 2 CLKINVX3 $T=1255980 2025520 1 0 $X=1255978 $Y=2020080
X1458 4598 4 3987 2 CLKINVX3 $T=1257300 2045680 1 0 $X=1257298 $Y=2040240
X1459 281 4 282 2 CLKINVX3 $T=1364880 2106160 0 0 $X=1364878 $Y=2105758
X1460 283 4 284 2 CLKINVX3 $T=1366200 2166640 0 0 $X=1366198 $Y=2166238
X1461 291 4 292 2 CLKINVX3 $T=1383360 2086000 1 0 $X=1383358 $Y=2080560
X1462 5082 4 195 2 CLKINVX3 $T=1428240 2086000 1 0 $X=1428238 $Y=2080560
X1463 244 4 263 2 CLKINVX3 $T=1440780 2035600 1 0 $X=1440778 $Y=2030160
X1464 4469 4 251 2 CLKINVX3 $T=1452660 2086000 1 0 $X=1452658 $Y=2080560
X1465 324 4 323 2 CLKINVX3 $T=1468500 2116240 0 0 $X=1468498 $Y=2115838
X1466 285 4 326 2 CLKINVX3 $T=1475100 2136400 0 0 $X=1475098 $Y=2135998
X1467 334 4 5493 2 CLKINVX3 $T=1489620 2116240 1 180 $X=1487640 $Y=2115838
X1468 370 4 311 2 CLKINVX3 $T=1581360 2005360 1 180 $X=1579380 $Y=2004958
X1469 6099 4 5573 2 CLKINVX3 $T=1584000 2186800 0 0 $X=1583998 $Y=2186398
X1470 374 4 382 2 CLKINVX3 $T=1599840 2065840 0 180 $X=1597860 $Y=2060400
X1471 373 4 6325 2 CLKINVX3 $T=1620960 2106160 0 0 $X=1620958 $Y=2105758
X1472 6415 4 378 2 CLKINVX3 $T=1658580 2186800 0 0 $X=1658578 $Y=2186398
X1473 407 4 293 2 CLKINVX3 $T=1683660 2217040 1 180 $X=1681680 $Y=2216638
X1474 6623 4 322 2 CLKINVX3 $T=1694220 2156560 0 0 $X=1694218 $Y=2156158
X1475 410 4 418 2 CLKINVX3 $T=1706100 2146480 0 0 $X=1706098 $Y=2146078
X1476 408 4 227 2 CLKINVX3 $T=1718640 2217040 1 0 $X=1718638 $Y=2211600
X1477 6836 4 310 2 CLKINVX3 $T=1724580 2206960 0 180 $X=1722600 $Y=2201520
X1478 6941 4 309 2 CLKINVX3 $T=1759560 2136400 0 0 $X=1759558 $Y=2135998
X1479 444 4 477 2 CLKINVX3 $T=1875060 2186800 1 0 $X=1875058 $Y=2181360
X1480 493 4 303 2 CLKINVX3 $T=1877040 2005360 0 180 $X=1875060 $Y=1999920
X1481 455 4 461 2 CLKINVX3 $T=1903440 2166640 1 0 $X=1903438 $Y=2161200
X1482 458 4 441 2 CLKINVX3 $T=1912680 2166640 0 0 $X=1912678 $Y=2166238
X1483 7775 4 7777 2 CLKINVX3 $T=1937760 2035600 0 0 $X=1937758 $Y=2035198
X1484 7732 4 7845 2 CLKINVX3 $T=1937760 2116240 1 0 $X=1937758 $Y=2110800
X1485 611 4 8670 2 CLKINVX3 $T=2143680 2065840 0 180 $X=2141700 $Y=2060400
X1486 9215 4 9230 2 CLKINVX3 $T=2214960 2146480 0 0 $X=2214958 $Y=2146078
X1487 9487 4 9655 2 CLKINVX3 $T=2295480 2217040 1 0 $X=2295478 $Y=2211600
X1488 9587 4 9542 2 CLKINVX3 $T=2296140 2005360 1 0 $X=2296138 $Y=1999920
X1489 663 4 668 2 CLKINVX3 $T=2374680 1995280 1 0 $X=2374678 $Y=1989840
X1490 10294 4 10442 2 CLKINVX3 $T=2463120 2126320 0 0 $X=2463118 $Y=2125918
X1491 2841 2839 4 2 2935 AND2X1 $T=924000 2106160 1 0 $X=923998 $Y=2100720
X1492 3880 3781 4 2 3968 AND2X1 $T=1120020 2075920 1 0 $X=1120018 $Y=2070480
X1493 125 3666 4 2 3961 AND2X1 $T=1130580 2196880 1 0 $X=1130578 $Y=2191440
X1494 131 3818 4 2 175 AND2X1 $T=1153680 2206960 1 180 $X=1151040 $Y=2206558
X1495 4696 4483 4 2 4742 AND2X1 $T=1286340 2015440 0 0 $X=1286338 $Y=2015038
X1496 251 252 4 2 4703 AND2X1 $T=1292940 2086000 0 180 $X=1290300 $Y=2080560
X1497 6480 6481 4 2 397 AND2X1 $T=1654620 2025520 1 0 $X=1654618 $Y=2020080
X1498 7614 499 4 2 7779 AND2X1 $T=1895520 2206960 0 0 $X=1895518 $Y=2206558
X1499 3414 3273 3420 4 123 2 AOI2BB1X4 $T=1017060 2206960 1 0 $X=1017058 $Y=2201520
X1500 2842 2829 4 2786 2828 2826 2 AOI22X1 $T=914760 2005360 1 180 $X=911460 $Y=2004958
X1501 5076 5040 4 4965 4998 5016 2 AOI22X1 $T=1353000 2075920 0 180 $X=1349700 $Y=2070480
X1502 369 334 4 301 366 5711 2 AOI22X1 $T=1571460 2106160 1 180 $X=1568160 $Y=2105758
X1503 392 394 4 395 262 6479 2 AOI22X1 $T=1650660 1995280 0 0 $X=1650658 $Y=1994878
X1504 393 394 4 395 233 6427 2 AOI22X1 $T=1650660 2005360 0 0 $X=1650658 $Y=2004958
X1505 6698 394 4 395 285 6620 2 AOI22X1 $T=1693560 2035600 0 180 $X=1690260 $Y=2030160
X1506 445 334 4 301 454 6835 2 AOI22X1 $T=1775400 2176720 1 180 $X=1772100 $Y=2176318
X1507 435 334 4 301 458 6857 2 AOI22X1 $T=1781340 2186800 0 0 $X=1781338 $Y=2186398
X1508 464 334 4 301 466 6757 2 AOI22X1 $T=1790580 2186800 0 0 $X=1790578 $Y=2186398
X1509 4683 4703 4719 4661 2 4 4758 OAI2BB2X1 $T=1286340 2096080 1 0 $X=1286338 $Y=2090640
X1510 8373 8352 8347 8393 2 4 8404 OAI2BB2X1 $T=2044680 2136400 1 0 $X=2044678 $Y=2130960
X1511 10975 10971 11004 10999 2 4 10978 OAI2BB2X1 $T=2562120 2055760 1 180 $X=2557500 $Y=2055358
X1512 608 567 639 9315 2 4 9336 ADDFXL $T=2226180 2075920 0 0 $X=2226178 $Y=2075518
X1513 164 166 2 4 4638 XNOR2XL $T=1259940 2217040 0 0 $X=1259938 $Y=2216638
X1514 251 4734 2 4 247 XNOR2XL $T=1288320 2005360 0 180 $X=1283040 $Y=1999920
X1515 413 6638 2 4 6617 XNOR2XL $T=1696860 2015440 0 180 $X=1691580 $Y=2010000
X1516 6761 6755 2 4 6770 XNOR2XL $T=1716000 2055760 0 0 $X=1715998 $Y=2055358
X1517 6760 6823 2 4 6711 XNOR2XL $T=1735800 2055760 1 180 $X=1730520 $Y=2055358
X1518 6925 6990 2 4 7026 XNOR2XL $T=1770120 2075920 0 0 $X=1770118 $Y=2075518
X1519 3140 264 4908 4 2 OR2X4 $T=1315380 2217040 1 0 $X=1315378 $Y=2211600
X1520 5260 7188 7170 4 2 OR2X4 $T=1804440 2126320 0 0 $X=1804438 $Y=2125918
X1521 498 500 7614 4 2 OR2X4 $T=1893540 2227120 1 0 $X=1893538 $Y=2221680
X1522 497 502 7607 4 2 OR2X4 $T=1898820 2126320 0 0 $X=1898818 $Y=2125918
X1523 507 510 7745 4 2 OR2X4 $T=1913340 2227120 0 0 $X=1913338 $Y=2226718
X1524 508 7746 7750 4 2 OR2X4 $T=1914660 2116240 1 0 $X=1914658 $Y=2110800
X1525 516 514 7810 4 2 OR2X4 $T=1933140 2055760 1 180 $X=1929180 $Y=2055358
X1526 520 517 7758 4 2 OR2X4 $T=1936440 2025520 1 180 $X=1932480 $Y=2025118
X1527 650 9489 9422 4 2 OR2X4 $T=2274360 2227120 1 180 $X=2270400 $Y=2226718
X1528 2524 2448 2444 2 4 100 OAI2BB1X4 $T=845460 2206960 0 180 $X=838860 $Y=2201520
X1529 8628 8474 8668 2 4 8677 OAI2BB1X4 $T=2098140 2035600 1 0 $X=2098138 $Y=2030160
X1530 615 9044 9039 2 4 9185 OAI2BB1X4 $T=2179320 2206960 0 0 $X=2179318 $Y=2206558
X1531 9230 9656 9657 2 4 9667 OAI2BB1X4 $T=2298780 2146480 0 0 $X=2298778 $Y=2146078
X1532 6326 347 2 4 INVX8 $T=1620960 2156560 0 0 $X=1620958 $Y=2156158
X1533 530 7851 2 4 INVX8 $T=1953600 2206960 0 0 $X=1953598 $Y=2206558
X1534 10395 688 2 4 INVX8 $T=2461140 2156560 1 0 $X=2461138 $Y=2151120
X1535 10317 10315 10297 685 4 2 MX2X4 $T=2443980 2176720 1 180 $X=2437380 $Y=2176318
X1536 2868 2863 106 2 4 NAND2BX2 $T=921360 2227120 0 180 $X=917400 $Y=2221680
X1537 3539 3543 3482 2 4 NAND2BX2 $T=1043460 2166640 1 0 $X=1043458 $Y=2161200
X1538 2845 2834 2832 2831 4 2 OAI2BB1X2 $T=916740 2096080 0 180 $X=912120 $Y=2090640
X1539 3118 3117 3108 115 4 2 OAI2BB1X2 $T=964260 2176720 1 180 $X=959640 $Y=2176318
X1540 3184 117 3109 3139 4 2 OAI2BB1X2 $T=976800 2186800 0 0 $X=976798 $Y=2186398
X1541 8407 8307 8437 8474 4 2 OAI2BB1X2 $T=2049960 2035600 0 0 $X=2049958 $Y=2035198
X1542 4505 233 231 2 4 4618 AND3X2 $T=1251360 2086000 0 0 $X=1251358 $Y=2085598
X1543 9020 9043 9098 2 4 9215 AND3X2 $T=2191860 2146480 1 0 $X=2191858 $Y=2141040
X1544 9654 9230 9494 2 4 9663 AND3X2 $T=2299440 2156560 0 0 $X=2299438 $Y=2156158
X1545 3818 131 2 4 4075 XOR2XL $T=1151040 2196880 0 0 $X=1151038 $Y=2196478
X1546 367 365 2 4 6058 XOR2XL $T=1570140 2227120 0 180 $X=1564860 $Y=2221680
X1547 6254 6299 2 4 385 XOR2XL $T=1618320 1995280 0 0 $X=1618318 $Y=1994878
X1548 6710 6717 2 4 6621 XOR2XL $T=1709400 2045680 1 180 $X=1704120 $Y=2045278
X1549 423 6758 2 4 6720 XOR2XL $T=1719960 2005360 0 180 $X=1714680 $Y=1999920
X1550 6828 6833 2 4 6768 XOR2XL $T=1738440 2075920 1 180 $X=1733160 $Y=2075518
X1551 540 8021 2 4 6807 XOR2XL $T=1974060 2005360 0 180 $X=1968780 $Y=1999920
X1552 8569 8571 2 4 8595 XOR2XL $T=2086260 2136400 0 0 $X=2086258 $Y=2135998
X1553 179 104 131 4170 4120 4 2 4109 SDFFRHQXL $T=1186680 2025520 0 180 $X=1170180 $Y=2020080
X1554 179 104 187 4175 4120 4 2 4087 SDFFRHQXL $T=1187340 2005360 1 180 $X=1170840 $Y=2004958
X1555 179 104 3666 4302 4120 4 2 4221 SDFFRHQXL $T=1211100 2055760 1 180 $X=1194600 $Y=2055358
X1556 179 104 186 4297 4120 4 2 4355 SDFFRHQXL $T=1199220 2106160 0 0 $X=1199218 $Y=2105758
X1557 179 104 149 4299 4120 4 2 4360 SDFFRHQXL $T=1199880 2096080 0 0 $X=1199878 $Y=2095678
X1558 239 104 5572 5556 4120 4 2 5469 SDFFRHQXL $T=1459260 2156560 1 180 $X=1442760 $Y=2156158
X1559 239 104 304 5489 4120 4 2 5594 SDFFRHQXL $T=1443420 2206960 1 0 $X=1443418 $Y=2201520
X1560 239 104 285 5689 4120 4 2 5778 SDFFRHQXL $T=1485000 2136400 0 0 $X=1484998 $Y=2135998
X1561 239 104 5082 5693 4120 4 2 5783 SDFFRHQXL $T=1486320 2086000 0 0 $X=1486318 $Y=2085598
X1562 239 104 233 5639 4120 4 2 5785 SDFFRHQXL $T=1487640 2156560 0 0 $X=1487638 $Y=2156158
X1563 239 104 262 5862 4120 4 2 5809 SDFFRHQXL $T=1527240 2136400 1 180 $X=1510740 $Y=2135998
X1564 239 104 353 5950 4120 4 2 6018 SDFFRHQXL $T=1538460 2136400 1 0 $X=1538458 $Y=2130960
X1565 239 104 386 6358 4120 4 2 6405 SDFFRHQXL $T=1626240 2146480 0 0 $X=1626238 $Y=2146078
X1566 239 104 6315 6359 4120 4 2 6389 SDFFRHQXL $T=1626900 2086000 0 0 $X=1626898 $Y=2085598
X1567 239 104 383 6269 4120 4 2 6515 SDFFRHQXL $T=1646040 2086000 1 0 $X=1646038 $Y=2080560
X1568 239 104 360 6579 4120 4 2 6633 SDFFRHQXL $T=1710060 2116240 1 180 $X=1693560 $Y=2115838
X1569 239 104 400 6712 4120 4 2 6623 SDFFRHQXL $T=1710060 2136400 0 180 $X=1693560 $Y=2130960
X1570 239 104 407 6713 4120 4 2 6635 SDFFRHQXL $T=1710720 2217040 1 180 $X=1694220 $Y=2216638
X1571 239 104 408 6724 4120 4 2 6616 SDFFRHQXL $T=1714020 2206960 1 180 $X=1697520 $Y=2206558
X1572 239 104 369 6756 4120 4 2 6851 SDFFRHQXL $T=1712040 2106160 0 0 $X=1712038 $Y=2105758
X1573 239 104 428 6803 4120 4 2 6746 SDFFRHQXL $T=1731180 2136400 1 180 $X=1714680 $Y=2135998
X1574 239 104 349 6864 4120 4 2 6941 SDFFRHQXL $T=1739760 2146480 1 0 $X=1739758 $Y=2141040
X1575 239 104 437 6888 4120 4 2 6988 SDFFRHQXL $T=1745040 2217040 0 0 $X=1745038 $Y=2216638
X1576 239 104 456 7075 4120 4 2 7019 SDFFRHQXL $T=1793880 2196880 1 180 $X=1777380 $Y=2196478
X1577 239 104 452 7217 4120 4 2 7273 SDFFRHQXL $T=1809720 2186800 1 0 $X=1809718 $Y=2181360
X1578 103 4 104 2 BUFX3 $T=872520 1995280 0 0 $X=872518 $Y=1994878
X1579 3666 4 135 2 BUFX3 $T=1069200 2055760 0 0 $X=1069198 $Y=2055358
X1580 183 4 4120 2 BUFX3 $T=1174140 2005360 1 0 $X=1174138 $Y=1999920
X1581 192 4 3937 2 BUFX3 $T=1191300 2015440 1 180 $X=1188660 $Y=2015038
X1582 186 4 3561 2 BUFX3 $T=1195920 2106160 0 0 $X=1195918 $Y=2105758
X1583 4221 4 125 2 BUFX3 $T=1197240 2065840 1 0 $X=1197238 $Y=2060400
X1584 4360 4 3666 2 BUFX3 $T=1202520 2086000 0 180 $X=1199880 $Y=2080560
X1585 300 4 252 2 BUFX3 $T=1390620 2065840 1 180 $X=1387980 $Y=2065438
X1586 5469 4 233 2 BUFX3 $T=1440780 2146480 1 180 $X=1438140 $Y=2146078
X1587 5575 4 4469 2 BUFX3 $T=1462560 2196880 0 0 $X=1462558 $Y=2196478
X1588 356 4 4196 2 BUFX3 $T=1537800 2156560 0 180 $X=1535160 $Y=2151120
X1589 5082 4 368 2 BUFX3 $T=1561560 2196880 1 0 $X=1561558 $Y=2191440
X1590 370 4 4209 2 BUFX3 $T=1582020 2025520 0 180 $X=1579380 $Y=2020080
X1591 6099 4 6345 2 BUFX3 $T=1619640 2186800 0 0 $X=1619638 $Y=2186398
X1592 6326 4 6338 2 BUFX3 $T=1624920 2156560 0 0 $X=1624918 $Y=2156158
X1593 6315 4 396 2 BUFX3 $T=1660560 2146480 1 0 $X=1660558 $Y=2141040
X1594 6415 4 6591 2 BUFX3 $T=1660560 2186800 0 0 $X=1660558 $Y=2186398
X1595 6616 4 407 2 BUFX3 $T=1689600 2206960 1 180 $X=1686960 $Y=2206558
X1596 395 4 6622 2 BUFX3 $T=1689600 2065840 1 0 $X=1689598 $Y=2060400
X1597 6635 4 337 2 BUFX3 $T=1693560 2227120 1 180 $X=1690920 $Y=2226718
X1598 6988 4 456 2 BUFX3 $T=1776060 2217040 0 0 $X=1776058 $Y=2216638
X1599 7019 4 462 2 BUFX3 $T=1783980 2217040 1 0 $X=1783978 $Y=2211600
X1600 7273 4 438 2 BUFX3 $T=1835460 2186800 1 0 $X=1835458 $Y=2181360
X1601 568 4 8456 2 BUFX3 $T=2058540 2075920 1 0 $X=2058538 $Y=2070480
X1602 601 4 8704 2 BUFX3 $T=2112000 2035600 0 180 $X=2109360 $Y=2030160
X1603 9454 4 7528 2 BUFX3 $T=2264460 2035600 1 180 $X=2261820 $Y=2035198
X1604 9909 4 7587 2 BUFX3 $T=2350920 2025520 0 180 $X=2348280 $Y=2020080
X1605 394 6711 4 363 409 6622 5082 6618 2 AOI222X2 $T=1698840 2055760 1 180 $X=1689600 $Y=2055358
X1606 304 4 335 5718 2 NOR2BXL $T=1490280 2217040 1 0 $X=1490278 $Y=2211600
X1607 5082 4 363 6033 2 NOR2BXL $T=1558920 2196880 1 0 $X=1558918 $Y=2191440
X1608 6099 4 233 6053 2 NOR2BXL $T=1575420 2176720 0 180 $X=1572780 $Y=2171280
X1609 3057 3058 2 4 2984 3108 AOI2BB1X1 $T=952380 2176720 0 0 $X=952378 $Y=2176318
X1610 3486 3508 2 4 3513 3549 AOI2BB1X1 $T=1037520 2005360 1 0 $X=1037518 $Y=1999920
X1611 3532 3389 2 4 3535 3658 AOI2BB1X1 $T=1041480 2065840 1 0 $X=1041478 $Y=2060400
X1612 5001 5027 2 4 5000 5099 AOI2BB1X1 $T=1346400 2196880 0 0 $X=1346398 $Y=2196478
X1613 347 262 2 4 5887 5894 AOI2BB1X1 $T=1527900 2166640 1 0 $X=1527898 $Y=2161200
X1614 351 6012 2 4 5867 5980 AOI2BB1X1 $T=1552980 2217040 1 180 $X=1549680 $Y=2216638
X1615 5493 312 2 5442 4 5399 5218 OAI211X1 $T=1434840 2116240 1 180 $X=1430880 $Y=2115838
X1616 5493 5508 2 5492 4 5490 5488 OAI211X1 $T=1447380 2116240 0 180 $X=1443420 $Y=2110800
X1617 5493 5509 2 5339 4 5487 5489 OAI211X1 $T=1447380 2176720 1 180 $X=1443420 $Y=2176318
X1618 5493 5573 2 5364 4 5555 5556 OAI211X1 $T=1455300 2176720 0 180 $X=1451340 $Y=2171280
X1619 5493 347 2 5324 4 5554 5639 OAI211X1 $T=1476420 2166640 0 180 $X=1472460 $Y=2161200
X1620 5493 5656 2 5363 4 5640 5618 OAI211X1 $T=1476420 2176720 1 180 $X=1472460 $Y=2176318
X1621 5493 343 2 5823 4 5819 5862 OAI211X1 $T=1511400 2116240 0 0 $X=1511398 $Y=2115838
X1622 2967 2885 93 2 4 3329 XNOR3X2 $T=955020 2005360 0 0 $X=955018 $Y=2004958
X1623 8373 8352 8347 2 4 8327 XNOR3X2 $T=2047320 2146480 0 180 $X=2035440 $Y=2141040
X1624 714 715 649 2 4 10922 XNOR3X2 $T=2535720 1995280 0 0 $X=2535718 $Y=1994878
X1625 11062 10975 10971 2 4 11021 XNOR3X2 $T=2574660 2055760 0 180 $X=2562780 $Y=2050320
X1626 11175 10844 11020 2 4 11163 XNOR3X2 $T=2608980 2055760 1 180 $X=2597100 $Y=2055358
X1627 312 4 300 262 347 5887 2 AOI22XL $T=1527900 2176720 1 0 $X=1527898 $Y=2171280
X1628 349 4 334 301 324 5941 2 AOI22XL $T=1535820 2116240 0 0 $X=1535818 $Y=2115838
X1629 364 4 6052 6052 4469 5934 2 AOI22XL $T=1564860 2166640 0 180 $X=1561560 $Y=2161200
X1630 383 4 334 301 374 6143 2 AOI22XL $T=1589280 2065840 1 180 $X=1585980 $Y=2065438
X1631 386 4 334 301 410 6478 2 AOI22XL $T=1695540 2146480 1 180 $X=1692240 $Y=2146078
X1632 438 4 334 301 444 6897 2 AOI22XL $T=1756260 2186800 0 180 $X=1752960 $Y=2181360
X1633 462 4 334 301 449 6834 2 AOI22XL $T=1768800 2186800 0 180 $X=1765500 $Y=2181360
X1634 452 4 334 301 451 6791 2 AOI22XL $T=1771440 2186800 1 180 $X=1768140 $Y=2186398
X1635 456 4 334 301 455 6882 2 AOI22XL $T=1778040 2166640 1 180 $X=1774740 $Y=2166238
X1636 4087 131 2 4 BUFX4 $T=1156980 2015440 0 180 $X=1153680 $Y=2010000
X1637 4109 138 2 4 BUFX4 $T=1162260 2025520 0 180 $X=1158960 $Y=2020080
X1638 4355 149 2 4 BUFX4 $T=1205160 2116240 1 180 $X=1201860 $Y=2115838
X1639 5594 276 2 4 BUFX4 $T=1450020 2227120 0 180 $X=1446720 $Y=2221680
X1640 5785 262 2 4 BUFX4 $T=1496220 2176720 1 180 $X=1492920 $Y=2176318
X1641 5809 285 2 4 BUFX4 $T=1511400 2146480 1 0 $X=1511398 $Y=2141040
X1642 6315 384 2 4 BUFX4 $T=1619640 2136400 1 0 $X=1619638 $Y=2130960
X1643 6515 363 2 4 BUFX4 $T=1671120 2086000 1 0 $X=1671118 $Y=2080560
X1644 6033 285 2 6033 343 5929 4 OAI22XL $T=1552320 2196880 0 180 $X=1548360 $Y=2191440
X1645 3987 2 130 4 CLKINVX8 $T=1143120 2015440 0 0 $X=1143118 $Y=2015038
X1646 5656 2 364 4 CLKINVX8 $T=1576740 2196880 1 0 $X=1576738 $Y=2191440
X1647 6315 2 312 4 CLKINVX8 $T=1609740 2136400 0 180 $X=1605780 $Y=2130960
X1648 399 396 300 395 401 394 403 2 4 AOI222X4 $T=1657920 1995280 1 0 $X=1657918 $Y=1989840
X1649 6164 399 251 395 404 394 405 2 4 AOI222X4 $T=1673100 1995280 1 0 $X=1673098 $Y=1989840
X1650 409 371 395 276 6617 394 411 2 4 AOI222X4 $T=1686960 2025520 1 0 $X=1686958 $Y=2020080
X1651 328 409 395 280 6621 394 427 2 4 AOI222X4 $T=1687620 2055760 1 0 $X=1687618 $Y=2050320
X1652 409 349 395 294 6931 394 446 2 4 AOI222X4 $T=1752960 2055760 0 0 $X=1752958 $Y=2055358
X1653 369 409 5953 395 6943 394 447 2 4 AOI222X4 $T=1755600 2045680 0 0 $X=1755598 $Y=2045278
X1654 445 409 314 395 6947 394 453 2 4 AOI222X4 $T=1756920 1995280 1 0 $X=1756918 $Y=1989840
X1655 386 409 311 395 6948 394 450 2 4 AOI222X4 $T=1756920 2005360 1 0 $X=1756918 $Y=1999920
X1656 383 409 295 395 6949 394 448 2 4 AOI222X4 $T=1756920 2015440 1 0 $X=1756918 $Y=2010000
X1657 239 104 325 6867 4120 11309 2 4 6836 SDFFRXL $T=1756920 2206960 0 180 $X=1738440 $Y=2201520
X1658 4196 193 191 2 182 4 194 196 4166 OAI222XL $T=1189980 2035600 0 0 $X=1189978 $Y=2035198
X1659 170 191 193 2 4209 4 197 196 4121 OAI222XL $T=1190640 2086000 0 0 $X=1190638 $Y=2085598
X1660 3794 191 193 2 195 4 200 196 4175 OAI222XL $T=1191960 2005360 1 0 $X=1191958 $Y=1999920
X1661 3765 191 193 2 4320 4 202 196 4299 OAI222XL $T=1203840 2086000 0 0 $X=1203838 $Y=2085598
X1662 231 193 191 2 137 4 205 196 4302 OAI222XL $T=1216380 2035600 1 180 $X=1211100 $Y=2035198
X1663 218 193 191 2 3638 4 210 196 4297 OAI222XL $T=1223640 2086000 1 180 $X=1218360 $Y=2085598
X1664 128 191 193 2 213 4 216 196 4154 OAI222XL $T=1220340 2075920 1 0 $X=1220338 $Y=2070480
X1665 150 191 193 2 215 4 217 196 4170 OAI222XL $T=1221000 2045680 1 0 $X=1220998 $Y=2040240
X1666 152 191 193 2 4469 4 222 196 219 OAI222XL $T=1229580 1995280 1 0 $X=1229578 $Y=1989840
X1667 227 193 191 2 3795 4 221 196 4411 OAI222XL $T=1236180 2045680 0 180 $X=1230900 $Y=2040240
X1668 244 193 191 2 4604 4 240 196 241 OAI222XL $T=1273140 2035600 1 180 $X=1267860 $Y=2035198
X1669 3987 191 193 2 255 4 258 196 4635 OAI222XL $T=1291620 2045680 1 0 $X=1291618 $Y=2040240
X1670 3958 191 193 2 268 4 269 196 4947 OAI222XL $T=1318680 2045680 1 0 $X=1318678 $Y=2040240
X1671 5800 276 5509 2 5800 4 5509 276 5799 OAI222XL $T=1510080 2206960 0 180 $X=1504800 $Y=2201520
X1672 5799 231 328 2 5799 4 231 328 5839 OAI222XL $T=1513380 2206960 0 0 $X=1513378 $Y=2206558
X1673 4196 5983 349 2 5983 4 4196 349 6012 OAI222XL $T=1552980 2196880 1 180 $X=1547700 $Y=2196478
X1674 6079 285 6079 2 343 4 343 285 5983 OAI222XL $T=1564860 2196880 1 180 $X=1559580 $Y=2196478
X1675 284 376 6216 2 5573 4 303 6248 6212 OAI222XL $T=1598520 2166640 0 0 $X=1598518 $Y=2166238
X1676 376 242 216 2 6248 4 6216 5509 6250 OAI222XL $T=1605120 2176720 1 180 $X=1599840 $Y=2176318
X1677 376 266 222 2 6255 4 6216 5656 6247 OAI222XL $T=1607760 2146480 1 180 $X=1602480 $Y=2146078
X1678 376 282 258 2 6256 4 6216 312 6258 OAI222XL $T=1608420 2106160 1 180 $X=1603140 $Y=2105758
X1679 376 292 200 2 6256 4 6215 5508 6269 OAI222XL $T=1611720 2086000 0 180 $X=1606440 $Y=2080560
X1680 382 376 6215 2 6287 4 217 6248 6277 OAI222XL $T=1614360 2065840 0 180 $X=1609080 $Y=2060400
X1681 376 257 269 2 6255 4 6216 347 6295 OAI222XL $T=1615680 2156560 1 180 $X=1610400 $Y=2156158
X1682 376 260 240 2 6256 4 6216 378 6296 OAI222XL $T=1616340 2166640 1 180 $X=1611060 $Y=2166238
X1683 376 234 205 2 6255 4 6325 6395 6359 OAI222XL $T=1634820 2106160 0 0 $X=1634818 $Y=2105758
X1684 376 398 202 2 6248 4 6325 343 6501 OAI222XL $T=1661220 2116240 1 0 $X=1661218 $Y=2110800
X1685 376 406 210 2 6256 4 6325 351 6579 OAI222XL $T=1683660 2116240 0 180 $X=1678380 $Y=2110800
X1686 376 323 194 2 6255 4 6325 433 6756 OAI222XL $T=1737120 2116240 1 0 $X=1737118 $Y=2110800
X1687 376 418 197 2 6248 4 6325 434 6803 OAI222XL $T=1737780 2146480 0 0 $X=1737778 $Y=2146078
X1688 376 441 431 2 6248 4 6325 443 6858 OAI222XL $T=1746360 2166640 0 0 $X=1746358 $Y=2166238
X1689 376 461 436 2 6256 4 6325 463 6888 OAI222XL $T=1782660 2166640 1 0 $X=1782658 $Y=2161200
X1690 376 467 429 2 6256 4 6325 468 7075 OAI222XL $T=1794540 2166640 1 0 $X=1794538 $Y=2161200
X1691 376 472 426 2 6255 4 6325 471 7191 OAI222XL $T=1809060 2176720 1 180 $X=1803780 $Y=2176318
X1692 376 475 421 2 6255 4 6325 480 7215 OAI222XL $T=1816980 2146480 0 0 $X=1816978 $Y=2146078
X1693 376 476 221 2 6256 4 6325 481 7213 OAI222XL $T=1816980 2166640 0 0 $X=1816978 $Y=2166238
X1694 376 477 439 2 6255 4 6325 482 7217 OAI222XL $T=1818300 2176720 0 0 $X=1818298 $Y=2176318
X1695 6427 6425 2 4 391 AND2X4 $T=1647360 2005360 0 0 $X=1647358 $Y=2004958
X1696 8718 8674 2 4 8742 AND2X4 $T=2110680 2217040 1 0 $X=2110678 $Y=2211600
X1697 8005 4 2 542 BUFX8 $T=1969440 2005360 0 0 $X=1969438 $Y=2004958
X1698 544 4 2 546 BUFX8 $T=1981320 2156560 1 0 $X=1981318 $Y=2151120
X1699 231 328 2 5858 4 5828 5841 OAI211XL $T=1519320 2196880 1 0 $X=1519318 $Y=2191440
X1700 239 104 4485 4635 4120 4 2 4598 SDFFRHQX1 $T=1267860 2055760 0 180 $X=1251360 $Y=2050320
X1701 179 104 182 4154 4120 3815 2 4 SDFFRHQX2 $T=1182060 2075920 0 180 $X=1162260 $Y=2070480
X1702 239 104 337 6858 4120 435 2 4 SDFFRHQX2 $T=1738440 2217040 1 0 $X=1738438 $Y=2211600
X1703 203 2421 2 4 BUFX12 $T=1208460 2015440 0 0 $X=1208458 $Y=2015038
X1704 179 3815 104 4121 4120 4 2 186 SDFFRHQX4 $T=1161600 2096080 0 0 $X=1161598 $Y=2095678
X1705 239 130 104 4947 4120 4 2 157 SDFFRHQX4 $T=1331880 2055760 0 180 $X=1307460 $Y=2050320
X1706 239 157 104 5218 4120 4 2 300 SDFFRHQX4 $T=1380720 2116240 0 0 $X=1380718 $Y=2115838
X1707 239 4469 104 5400 4120 4 2 280 SDFFRHQX4 $T=1431540 2196880 1 180 $X=1407120 $Y=2196478
X1708 239 280 104 5406 4120 4 2 304 SDFFRHQX4 $T=1431540 2206960 0 180 $X=1407120 $Y=2201520
X1709 239 300 104 5488 4120 4 2 5082 SDFFRHQX4 $T=1461900 2136400 1 180 $X=1437480 $Y=2135998
X1710 239 294 104 6247 4120 4 2 6164 SDFFRHQX4 $T=1611060 2126320 1 180 $X=1586640 $Y=2125918
X1711 239 311 104 6212 4120 4 2 6099 SDFFRHQX4 $T=1595220 2186800 0 0 $X=1595218 $Y=2186398
X1712 239 6415 104 6295 4120 4 2 6326 SDFFRHQX4 $T=1646700 2176720 1 180 $X=1622280 $Y=2176318
X1713 239 6164 104 6258 4120 4 2 6315 SDFFRHQX4 $T=1623600 2126320 0 0 $X=1623598 $Y=2125918
X1714 239 6345 104 6296 4120 4 2 6415 SDFFRHQX4 $T=1626900 2186800 0 0 $X=1626898 $Y=2186398
X1715 239 328 104 6277 4120 4 2 383 SDFFRHQX4 $T=1627560 2065840 1 0 $X=1627558 $Y=2060400
X1716 239 363 104 6501 4120 4 2 400 SDFFRHQX4 $T=1655940 2136400 1 0 $X=1655938 $Y=2130960
X1717 239 6326 104 6250 4120 4 2 371 SDFFRHQX4 $T=1659900 2186800 1 0 $X=1659898 $Y=2181360
X1718 239 371 104 6695 4120 4 2 408 SDFFRHQX4 $T=1706100 2186800 1 180 $X=1681680 $Y=2186398
X1719 239 435 104 6860 4120 4 2 325 SDFFRHQX4 $T=1739100 2196880 0 0 $X=1739098 $Y=2196478
X1720 239 445 104 7191 4120 4 2 452 SDFFRHQX4 $T=1806420 2196880 1 0 $X=1806418 $Y=2191440
X1721 239 462 104 7213 4120 4 2 445 SDFFRHQX4 $T=1807080 2196880 0 0 $X=1807078 $Y=2196478
X1722 239 438 104 7215 4120 4 2 464 SDFFRHQX4 $T=1808400 2156560 0 0 $X=1808398 $Y=2156158
X1723 269 5321 256 4 301 5324 2 AOI2BB2XL $T=1401180 2156560 0 0 $X=1401178 $Y=2156158
X1724 303 5321 283 4 301 5364 2 AOI2BB2XL $T=1409100 2166640 0 0 $X=1409098 $Y=2166238
X1725 5321 222 2 265 301 5363 4 AOI2BB2X2 $T=1406460 2156560 1 0 $X=1406458 $Y=2151120
X1726 8969 537 603 4 2 9095 ADDHX1 $T=2178660 2086000 1 0 $X=2178658 $Y=2080560
X1727 5272 294 280 227 268 288 5185 2 4 5123 CMPR42X1 $T=1396560 2045680 1 180 $X=1374120 $Y=2045278
X1728 5190 5209 289 5082 293 296 5272 2 4 298 CMPR42X1 $T=1378080 2025520 1 0 $X=1378078 $Y=2020080
X1729 5382 4469 297 295 5229 290 5190 2 4 287 CMPR42X1 $T=1400520 2005360 0 180 $X=1378080 $Y=1999920
X1730 5402 262 311 5383 5382 305 5361 2 4 302 CMPR42X1 $T=1430880 2005360 1 180 $X=1408440 $Y=2004958
X1731 315 5209 314 5459 5395 307 5402 2 4 306 CMPR42X1 $T=1442760 2015440 0 180 $X=1420320 $Y=2010000
X1732 5657 326 314 5616 5597 320 319 2 4 317 CMPR42X1 $T=1479720 2015440 1 180 $X=1457280 $Y=2015038
X1733 5595 321 5615 4196 5638 327 5657 2 4 330 CMPR42X1 $T=1461240 2035600 0 0 $X=1461238 $Y=2035198
X1734 5784 5082 5780 218 5690 331 5595 2 4 329 CMPR42X1 $T=1503480 2045680 1 180 $X=1481040 $Y=2045278
X1735 5801 5840 285 215 340 339 5784 2 4 336 CMPR42X1 $T=1522620 2015440 0 180 $X=1500180 $Y=2010000
X1736 5940 311 346 294 344 341 5801 2 4 338 CMPR42X1 $T=1527900 2005360 0 180 $X=1505460 $Y=1999920
X1737 362 360 321 295 227 355 5937 2 4 350 CMPR42X1 $T=1560240 1995280 0 180 $X=1537800 $Y=1989840
X1738 5937 314 337 5953 4209 357 5940 2 4 352 CMPR42X1 $T=1561560 2005360 1 180 $X=1539120 $Y=2004958
X1739 8614 584 567 565 8704 8719 8726 2 4 8692 CMPR42X1 $T=2095500 2096080 0 0 $X=2095498 $Y=2095678
X1740 8726 566 8456 603 583 8672 8669 2 4 8591 CMPR42X1 $T=2119260 2086000 1 180 $X=2096820 $Y=2085598
X1741 8924 583 8670 538 8804 8808 8614 2 4 8763 CMPR42X1 $T=2150280 2106160 0 180 $X=2127840 $Y=2100720
X1742 8973 8969 566 8852 8924 8892 8881 2 4 8829 CMPR42X1 $T=2167440 2086000 1 180 $X=2145000 $Y=2085598
X1743 9186 8670 8456 565 8997 8990 8974 2 4 8929 CMPR42X1 $T=2185920 2106160 0 180 $X=2163480 $Y=2100720
X1744 9212 626 567 8704 9095 9079 8973 2 4 8974 CMPR42X1 $T=2206380 2065840 1 180 $X=2183940 $Y=2065438
X1745 9081 9096 8704 9165 9167 9184 9189 2 4 9105 CMPR42X1 $T=2189220 2106160 0 0 $X=2189218 $Y=2105758
X1746 9096 583 567 538 8969 9167 9212 2 4 9164 CMPR42X1 $T=2193840 2086000 0 0 $X=2193838 $Y=2085598
X1747 9274 634 608 9186 9079 9166 9164 2 4 9035 CMPR42X1 $T=2219580 2096080 1 180 $X=2197140 $Y=2095678
X1748 9475 9336 9345 9081 9294 9280 9256 2 4 9253 CMPR42X1 $T=2246640 2116240 0 180 $X=2224200 $Y=2110800
X1749 9334 8670 566 565 626 9283 9183 2 4 9256 CMPR42X1 $T=2247300 2065840 1 180 $X=2224860 $Y=2065438
X1750 9345 622 566 538 9095 9294 9274 2 4 9189 CMPR42X1 $T=2247960 2106160 0 180 $X=2225520 $Y=2100720
X1751 9279 583 634 538 9334 9347 9315 2 4 9447 CMPR42X1 $T=2228820 2086000 0 0 $X=2228818 $Y=2085598
X1752 9530 9513 565 9475 9283 9455 9447 2 4 9360 CMPR42X1 $T=2281620 2106160 1 180 $X=2259180 $Y=2105758
X1753 9446 9456 9450 9347 9496 9514 9530 2 4 9508 CMPR42X1 $T=2261160 2116240 0 0 $X=2261158 $Y=2115838
X1754 9706 583 584 628 8704 9607 9279 2 4 9496 CMPR42X1 $T=2315280 2106160 0 180 $X=2292840 $Y=2100720
X1755 9721 584 634 656 8670 9608 9599 2 4 9580 CMPR42X1 $T=2315940 2075920 1 180 $X=2293500 $Y=2075518
X1756 9883 9520 9706 9607 9580 9661 9446 2 4 9600 CMPR42X1 $T=2319240 2116240 0 180 $X=2296800 $Y=2110800
X1757 9787 622 583 9608 9794 9873 9883 2 4 9809 CMPR42X1 $T=2330460 2106160 1 0 $X=2330458 $Y=2100720
X1758 9919 628 8670 9821 9721 9822 9521 2 4 9794 CMPR42X1 $T=2353560 2075920 0 180 $X=2331120 $Y=2070480
X1759 9991 8704 584 9976 9912 9932 9919 2 4 9913 CMPR42X1 $T=2375340 2045680 1 180 $X=2352900 $Y=2045278
X1760 10040 639 626 9822 9913 9935 9787 2 4 9861 CMPR42X1 $T=2376000 2086000 0 180 $X=2353560 $Y=2080560
X1761 9960 8670 656 9932 9977 10035 10040 2 4 10033 CMPR42X1 $T=2366100 2065840 0 0 $X=2366098 $Y=2065438
X1762 10144 8704 634 10046 10013 9998 9991 2 4 9977 CMPR42X1 $T=2391840 2055760 0 180 $X=2369400 $Y=2050320
X1763 10204 603 608 10135 9998 10054 9960 2 4 10036 CMPR42X1 $T=2405040 2075920 0 180 $X=2382600 $Y=2070480
X1764 10224 622 649 628 10160 10161 10144 2 4 10135 CMPR42X1 $T=2422860 2065840 0 180 $X=2400420 $Y=2060400
X1765 10296 10224 10274 10251 10161 10225 10204 2 4 10201 CMPR42X1 $T=2439360 2096080 0 180 $X=2416920 $Y=2090640
X1766 10438 10410 634 10391 10138 10314 10296 2 4 10290 CMPR42X1 $T=2459160 2086000 1 180 $X=2436720 $Y=2085598
X1767 10319 628 622 10393 10392 10418 10438 2 4 10435 CMPR42X1 $T=2442660 2075920 0 0 $X=2442658 $Y=2075518
X1768 10485 628 626 10473 10274 10554 10319 2 4 10518 CMPR42X1 $T=2470380 2086000 1 0 $X=2470378 $Y=2080560
X1769 10680 634 647 639 10410 10787 10485 2 4 10937 CMPR42X1 $T=2507340 2086000 1 0 $X=2507338 $Y=2080560
X1770 332 5808 2 4 CLKBUFX4 $T=1497540 2106160 1 0 $X=1497538 $Y=2100720
X1771 93 87 86 4 2 2073 ADDHX2 $T=830940 2015440 0 180 $X=819060 $Y=2010000
X1772 179 104 138 4166 4120 182 4 2 3818 SDFFRX1 $T=1184040 2055760 1 180 $X=1165560 $Y=2055358
X1773 179 104 125 4411 4120 3795 4 2 4485 SDFFRX1 $T=1220340 2055760 1 0 $X=1220338 $Y=2050320
X1774 239 104 295 5618 4120 5575 4 2 316 SDFFRX1 $T=1473120 2217040 0 180 $X=1454640 $Y=2211600
X1775 6285 312 5573 5656 4 2 377 NAND4BX4 $T=1603140 2196880 0 180 $X=1591260 $Y=2191440
.ENDS
***************************************
.SUBCKT XOR3X4 A B C Y VSS VDD
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57 2 4 29 30 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47
+ 48 49 50 51 52 54 56 60 61 62 65 66 67 68 69 72 73 74 78 80
+ 81 82 83 86 87 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106
+ 107 108 109 110 111 112 113 114 115 116 117 119 120 122 123 124 125 127 128 130
+ 131 132 133 134 136 137 140 143 144 145 147 148 149 152 153 154 155 157 158 159
+ 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 222 223 224 225 226 227 228 229 231 232 233 234 237 238 239 240 241 242 244 245
+ 246 248 250 251 252 254 255 256 257 258 260 261 265 267 268 269 270 271 272 273
+ 274 275 277 278 279 281 284 285 286 287 288 289 290 291 292 293 295 296 297 298
+ 299 300 301 302 303 304 305 306 307 308 309 310 311 313 314 316 317 319 320 321
+ 322 323 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 347 348 349 350 351 354 355 356 358 359 360 361 362 363 364 365 366
+ 367 368 369 370 372 373 374 375 376 377 378 379 380 381 382 383 387 388 390 391
+ 392 393 394 395 396 397 398 399 401 402 403 405 407 409 410 414 416 418 420 421
+ 423 424 425 426 427 428 430 431 432 433 434 435 436 437 438 439 440 441 442 443
+ 444 445 446 447 448 450 454 459 460 461 462 464 467 468 469 470 472 475 477 478
+ 479 482 484 485 489 490 493 494 495 498 501 502 503 505 506 507 511 514 519 525
+ 1414 1415
** N=28216 EP=382 IP=10170 FDC=0
X0 1559 4 1543 2 1558 NAND2X1 $T=702240 2297680 1 180 $X=700260 $Y=2297278
X1 1610 4 32 2 1572 NAND2X1 $T=712800 2297680 0 180 $X=710820 $Y=2292240
X2 1572 4 1625 2 1626 NAND2X1 $T=729300 2327920 0 0 $X=729298 $Y=2327518
X3 1625 4 1641 2 1642 NAND2X1 $T=734580 2327920 0 0 $X=734578 $Y=2327518
X4 1574 4 1657 2 1669 NAND2X1 $T=741180 2307760 0 0 $X=741178 $Y=2307358
X5 1736 4 1673 2 1684 NAND2X1 $T=752400 2297680 0 180 $X=750420 $Y=2292240
X6 1737 4 1638 2 1797 NAND2X1 $T=762960 2317840 1 0 $X=762958 $Y=2312400
X7 1724 4 1641 2 1759 NAND2X1 $T=762960 2338000 0 0 $X=762958 $Y=2337598
X8 1638 4 1641 2 1787 NAND2X1 $T=768240 2338000 1 0 $X=768238 $Y=2332560
X9 1785 4 1783 2 1825 NAND2X1 $T=786720 2297680 0 0 $X=786718 $Y=2297278
X10 2076 4 1738 2 2088 NAND2X1 $T=863940 2327920 0 0 $X=863938 $Y=2327518
X11 2059 4 2089 2 2107 NAND2X1 $T=866580 2307760 0 0 $X=866578 $Y=2307358
X12 2168 4 2104 2 2145 NAND2X1 $T=887040 2307760 0 180 $X=885060 $Y=2302320
X13 2176 4 2174 2 2179 NAND2X1 $T=896280 2338000 1 180 $X=894300 $Y=2337598
X14 2224 4 65 2 2259 NAND2X1 $T=911460 2247280 0 180 $X=909480 $Y=2241840
X15 2259 4 2228 2 2293 NAND2X1 $T=916080 2257360 1 0 $X=916078 $Y=2251920
X16 2296 4 2172 2 2309 NAND2X1 $T=926640 2317840 0 0 $X=926638 $Y=2317438
X17 2353 4 2355 2 2364 NAND2X1 $T=941160 2358160 0 0 $X=941158 $Y=2357758
X18 2352 4 2350 2 2380 NAND2X1 $T=946440 2327920 1 0 $X=946438 $Y=2322480
X19 2356 4 2353 2 2277 NAND2X1 $T=951720 2327920 0 0 $X=951718 $Y=2327518
X20 93 4 92 2 2652 NAND2X1 $T=1016400 2247280 0 180 $X=1014420 $Y=2241840
X21 2671 4 1874 2 2691 NAND2X1 $T=1024980 2368240 0 0 $X=1024978 $Y=2367838
X22 2691 4 2693 2 2669 NAND2X1 $T=1027620 2398480 1 0 $X=1027618 $Y=2393040
X23 2699 4 2697 2 2755 NAND2X1 $T=1032240 2297680 0 180 $X=1030260 $Y=2292240
X24 2716 4 2718 2 2692 NAND2X1 $T=1032240 2338000 0 0 $X=1032238 $Y=2337598
X25 2747 4 2734 2 2723 NAND2X1 $T=1040160 2388400 0 180 $X=1038180 $Y=2382960
X26 2733 4 2080 2 2747 NAND2X1 $T=1039500 2358160 0 0 $X=1039498 $Y=2357758
X27 2674 4 2690 2 2716 NAND2X1 $T=1040160 2327920 1 0 $X=1040158 $Y=2322480
X28 2807 4 1913 2 2769 NAND2X1 $T=1049400 2317840 1 180 $X=1047420 $Y=2317438
X29 2747 4 2770 2 2840 NAND2X1 $T=1048080 2378320 1 0 $X=1048078 $Y=2372880
X30 96 4 2765 2 2713 NAND2X1 $T=1053360 2257360 1 0 $X=1053358 $Y=2251920
X31 2866 4 2809 2 2672 NAND2X1 $T=1069200 2277520 1 0 $X=1069198 $Y=2272080
X32 2906 4 1902 2 2907 NAND2X1 $T=1079100 2398480 0 180 $X=1077120 $Y=2393040
X33 2904 4 1815 2 3004 NAND2X1 $T=1082400 2358160 1 0 $X=1082398 $Y=2352720
X34 2918 4 2922 2 2842 NAND2X1 $T=1083060 2277520 0 0 $X=1083058 $Y=2277118
X35 103 4 2937 2 2920 NAND2X1 $T=1087020 2267440 0 0 $X=1087018 $Y=2267038
X36 3004 4 3006 2 3046 NAND2X1 $T=1103520 2358160 1 0 $X=1103518 $Y=2352720
X37 2974 4 3020 2 3022 NAND2X1 $T=1107480 2297680 1 0 $X=1107478 $Y=2292240
X38 114 4 115 2 2997 NAND2X1 $T=1111440 2267440 1 0 $X=1111438 $Y=2262000
X39 2998 4 3038 2 3077 NAND2X1 $T=1112100 2348080 0 0 $X=1112098 $Y=2347678
X40 119 4 3083 2 3081 NAND2X1 $T=1127940 2247280 1 180 $X=1125960 $Y=2246878
X41 3126 4 120 2 3152 NAND2X1 $T=1153020 2267440 1 0 $X=1153018 $Y=2262000
X42 3220 4 3218 2 3219 NAND2X1 $T=1157640 2287600 0 180 $X=1155660 $Y=2282160
X43 3218 4 3224 2 3225 NAND2X1 $T=1160280 2307760 0 180 $X=1158300 $Y=2302320
X44 3258 4 3224 2 3270 NAND2X1 $T=1165560 2307760 0 180 $X=1163580 $Y=2302320
X45 133 4 130 2 3310 NAND2X1 $T=1182060 2257360 1 0 $X=1182058 $Y=2251920
X46 3308 4 2596 2 3311 NAND2X1 $T=1182060 2348080 0 0 $X=1182058 $Y=2347678
X47 136 4 137 2 3336 NAND2X1 $T=1189980 2257360 0 0 $X=1189978 $Y=2256958
X48 3425 4 3333 2 3426 NAND2X1 $T=1203840 2388400 0 0 $X=1203838 $Y=2387998
X49 3432 4 3299 2 3427 NAND2X1 $T=1205820 2297680 0 180 $X=1203840 $Y=2292240
X50 3442 4 3427 2 3445 NAND2X1 $T=1207140 2307760 0 180 $X=1205160 $Y=2302320
X51 3445 4 2191 2 3444 NAND2X1 $T=1209780 2368240 1 180 $X=1207800 $Y=2367838
X52 3450 4 3475 2 3442 NAND2X1 $T=1211760 2297680 0 0 $X=1211758 $Y=2297278
X53 144 4 145 2 3471 NAND2X1 $T=1215720 2247280 0 0 $X=1215718 $Y=2246878
X54 3497 4 2226 2 3495 NAND2X1 $T=1218360 2358160 0 180 $X=1216380 $Y=2352720
X55 3444 4 3425 2 3546 NAND2X1 $T=1217040 2388400 1 0 $X=1217038 $Y=2382960
X56 154 4 152 2 3593 NAND2X1 $T=1233540 2247280 1 180 $X=1231560 $Y=2246878
X57 3597 4 2445 2 3620 NAND2X1 $T=1241460 2348080 0 180 $X=1239480 $Y=2342640
X58 3593 4 3594 2 3619 NAND2X1 $T=1242120 2287600 1 0 $X=1242118 $Y=2282160
X59 3640 4 2597 2 3641 NAND2X1 $T=1248060 2368240 1 180 $X=1246080 $Y=2367838
X60 3627 4 3672 2 3741 NAND2X1 $T=1254000 2247280 1 0 $X=1253998 $Y=2241840
X61 159 4 158 2 3666 NAND2X1 $T=1255320 2257360 0 0 $X=1255318 $Y=2256958
X62 3684 4 3695 2 161 NAND2X1 $T=1259280 2388400 0 0 $X=1259278 $Y=2387998
X63 3526 4 3743 2 3742 NAND2X1 $T=1272480 2257360 1 180 $X=1270500 $Y=2256958
X64 3744 4 2366 2 3764 NAND2X1 $T=1277100 2348080 1 180 $X=1275120 $Y=2347678
X65 3728 4 3752 2 167 NAND2X1 $T=1275780 2408560 1 0 $X=1275778 $Y=2403120
X66 3695 4 3752 2 3801 NAND2X1 $T=1283700 2398480 0 0 $X=1283698 $Y=2398078
X67 3788 4 3752 2 171 NAND2X1 $T=1286340 2408560 1 0 $X=1286338 $Y=2403120
X68 2504 4 176 2 3897 NAND2X1 $T=1309440 2327920 1 180 $X=1307460 $Y=2327518
X69 2595 4 178 2 3972 NAND2X1 $T=1329900 2348080 0 0 $X=1329898 $Y=2347678
X70 3897 4 3961 2 3985 NAND2X1 $T=1338480 2317840 1 0 $X=1338478 $Y=2312400
X71 182 4 2328 2 4013 NAND2X1 $T=1345080 2307760 0 180 $X=1343100 $Y=2302320
X72 187 4 2455 2 4085 NAND2X1 $T=1357620 2297680 0 180 $X=1355640 $Y=2292240
X73 4165 4 4163 2 4007 NAND2X1 $T=1379400 2388400 1 0 $X=1379398 $Y=2382960
X74 4013 4 4066 2 4162 NAND2X1 $T=1380720 2297680 0 0 $X=1380718 $Y=2297278
X75 4183 4 4180 2 4082 NAND2X1 $T=1385340 2368240 0 180 $X=1383360 $Y=2362800
X76 4208 4 4229 2 202 NAND2X1 $T=1396560 2237200 0 0 $X=1396558 $Y=2236798
X77 4279 4 4274 2 4235 NAND2X1 $T=1402500 2388400 0 180 $X=1400520 $Y=2382960
X78 206 4 4278 2 4279 NAND2X1 $T=1404480 2358160 0 180 $X=1402500 $Y=2352720
X79 4292 4 4294 2 4210 NAND2X1 $T=1407120 2267440 0 0 $X=1407118 $Y=2267038
X80 4274 4 4305 2 4306 NAND2X1 $T=1409100 2378320 0 0 $X=1409098 $Y=2377918
X81 4318 4 4328 2 4330 NAND2X1 $T=1417680 2338000 0 0 $X=1417678 $Y=2337598
X82 4382 4 197 2 4208 NAND2X1 $T=1433520 2257360 0 0 $X=1433518 $Y=2256958
X83 4379 4 4363 2 4385 NAND2X1 $T=1435500 2348080 0 0 $X=1435498 $Y=2347678
X84 4464 4 4462 2 223 NAND2X1 $T=1454640 2408560 0 180 $X=1452660 $Y=2403120
X85 4538 4 232 2 4533 NAND2X1 $T=1479060 2388400 0 180 $X=1477080 $Y=2382960
X86 233 4 95 2 4538 NAND2X1 $T=1479060 2408560 0 0 $X=1479058 $Y=2408158
X87 4645 4 212 2 4642 NAND2X1 $T=1506780 2257360 1 180 $X=1504800 $Y=2256958
X88 4656 4 4660 2 4658 NAND2X1 $T=1510080 2378320 1 0 $X=1510078 $Y=2372880
X89 4678 4 4676 2 4657 NAND2X1 $T=1513380 2307760 1 180 $X=1511400 $Y=2307358
X90 4729 4 204 2 250 NAND2X1 $T=1527900 2247280 0 180 $X=1525920 $Y=2241840
X91 4745 4 4766 2 4706 NAND2X1 $T=1537800 2307760 1 0 $X=1537798 $Y=2302320
X92 4767 4 4769 2 4688 NAND2X1 $T=1538460 2388400 0 0 $X=1538458 $Y=2387998
X93 4777 4 4781 2 4656 NAND2X1 $T=1540440 2378320 1 0 $X=1540438 $Y=2372880
X94 4794 4 4789 2 4745 NAND2X1 $T=1545060 2307760 0 0 $X=1545058 $Y=2307358
X95 4854 4 4851 2 4714 NAND2X1 $T=1553640 2327920 1 0 $X=1553638 $Y=2322480
X96 4882 4 4824 2 4793 NAND2X1 $T=1563540 2277520 0 0 $X=1563538 $Y=2277118
X97 4902 4 4886 2 4852 NAND2X1 $T=1569480 2247280 1 180 $X=1567500 $Y=2246878
X98 4952 4 4901 2 4880 NAND2X1 $T=1579380 2237200 1 0 $X=1579378 $Y=2231760
X99 5033 4 5030 2 285 NAND2X1 $T=1605120 2247280 0 180 $X=1603140 $Y=2241840
X100 279 4 5032 2 5033 NAND2X1 $T=1605120 2257360 1 0 $X=1605118 $Y=2251920
X101 4708 4 5048 2 5046 NAND2X1 $T=1609740 2358160 0 0 $X=1609738 $Y=2357758
X102 279 4 281 2 5105 NAND2X1 $T=1626900 2277520 0 0 $X=1626898 $Y=2277118
X103 5098 4 5118 2 304 NAND2X1 $T=1629540 2368240 0 180 $X=1627560 $Y=2362800
X104 5068 4 5096 2 5098 NAND2X1 $T=1628880 2348080 0 0 $X=1628878 $Y=2347678
X105 270 4 5247 2 5263 NAND2X1 $T=1663200 2267440 1 0 $X=1663198 $Y=2262000
X106 304 4 302 2 5278 NAND2X1 $T=1668480 2398480 1 0 $X=1668478 $Y=2393040
X107 5069 4 5229 2 306 NAND2X1 $T=1671120 2398480 0 0 $X=1671118 $Y=2398078
X108 5426 4 5395 2 5328 NAND2X1 $T=1706760 2398480 0 180 $X=1704780 $Y=2393040
X109 5406 4 5323 2 5404 NAND2X1 $T=1708080 2348080 0 180 $X=1706100 $Y=2342640
X110 5519 4 5523 2 5504 NAND2X1 $T=1741080 2378320 0 180 $X=1739100 $Y=2372880
X111 5524 4 5422 2 5481 NAND2X1 $T=1741740 2398480 0 0 $X=1741738 $Y=2398078
X112 5601 4 5546 2 5676 NAND2X1 $T=1766160 2338000 0 0 $X=1766158 $Y=2337598
X113 278 4 5671 2 5658 NAND2X1 $T=1772760 2388400 0 0 $X=1772758 $Y=2387998
X114 5754 4 5847 2 5908 NAND2X1 $T=1815000 2317840 0 0 $X=1814998 $Y=2317438
X115 5847 4 5858 2 5862 NAND2X1 $T=1816980 2338000 1 0 $X=1816978 $Y=2332560
X116 351 4 3221 2 5927 NAND2X1 $T=1825560 2297680 0 0 $X=1825558 $Y=2297278
X117 6034 4 5863 2 6028 NAND2X1 $T=1859220 2348080 0 0 $X=1859218 $Y=2347678
X118 5833 4 5931 2 6015 NAND2X1 $T=1859220 2388400 0 0 $X=1859218 $Y=2387998
X119 360 4 3256 2 6061 NAND2X1 $T=1868460 2317840 0 0 $X=1868458 $Y=2317438
X120 5986 4 5830 2 6075 NAND2X1 $T=1872420 2398480 0 0 $X=1872418 $Y=2398078
X121 6061 4 6044 2 6057 NAND2X1 $T=1873740 2307760 0 0 $X=1873738 $Y=2307358
X122 6045 4 5910 2 6108 NAND2X1 $T=1876380 2338000 1 0 $X=1876378 $Y=2332560
X123 368 4 169 2 367 NAND2X1 $T=1892220 2237200 0 180 $X=1890240 $Y=2231760
X124 6116 4 6142 2 6202 NAND2X1 $T=1903440 2378320 1 0 $X=1903438 $Y=2372880
X125 373 4 190 2 372 NAND2X1 $T=1914660 2247280 0 180 $X=1912680 $Y=2241840
X126 6254 4 6260 2 6259 NAND2X1 $T=1921920 2307760 1 0 $X=1921918 $Y=2302320
X127 6191 4 6189 2 6285 NAND2X1 $T=1929840 2287600 1 0 $X=1929838 $Y=2282160
X128 6304 4 4065 2 6409 NAND2X1 $T=1957560 2277520 1 0 $X=1957558 $Y=2272080
X129 6410 4 3944 2 6449 NAND2X1 $T=1959540 2247280 0 0 $X=1959538 $Y=2246878
X130 6443 4 3931 2 6474 NAND2X1 $T=1970100 2368240 1 180 $X=1968120 $Y=2367838
X131 6474 4 6444 2 6486 NAND2X1 $T=1976700 2338000 1 180 $X=1974720 $Y=2337598
X132 398 4 3669 2 6534 NAND2X1 $T=1992540 2358160 1 0 $X=1992538 $Y=2352720
X133 6787 4 6802 2 6854 NAND2X1 $T=2077680 2297680 0 0 $X=2077678 $Y=2297278
X134 6857 4 6864 2 6885 NAND2X1 $T=2086920 2307760 0 0 $X=2086918 $Y=2307358
X135 6867 4 6866 2 6958 NAND2X1 $T=2088900 2358160 1 180 $X=2086920 $Y=2357758
X136 6804 4 6870 2 6858 NAND2X1 $T=2089560 2338000 1 0 $X=2089558 $Y=2332560
X137 6958 4 6948 2 6949 NAND2X1 $T=2104740 2358160 1 0 $X=2104738 $Y=2352720
X138 423 4 6959 2 428 NAND2X1 $T=2112660 2237200 1 0 $X=2112658 $Y=2231760
X139 6980 4 6947 2 7007 NAND2X1 $T=2119260 2277520 1 0 $X=2119258 $Y=2272080
X140 7006 4 7011 2 432 NAND2X1 $T=2123220 2408560 0 0 $X=2123218 $Y=2408158
X141 430 4 6994 2 7048 NAND2X1 $T=2131140 2247280 0 0 $X=2131138 $Y=2246878
X142 436 4 438 2 7088 NAND2X1 $T=2148960 2267440 1 0 $X=2148958 $Y=2262000
X143 7071 4 7138 2 440 NAND2X1 $T=2162820 2408560 1 180 $X=2160840 $Y=2408158
X144 7185 4 7167 2 7166 NAND2X1 $T=2175360 2287600 0 180 $X=2173380 $Y=2282160
X145 7166 4 7202 2 7203 NAND2X1 $T=2183280 2267440 1 0 $X=2183278 $Y=2262000
X146 7202 4 7284 2 7286 NAND2X1 $T=2205720 2267440 1 0 $X=2205718 $Y=2262000
X147 7303 4 7284 2 7283 NAND2X1 $T=2211660 2267440 1 180 $X=2209680 $Y=2267038
X148 7305 4 7315 2 7303 NAND2X1 $T=2220240 2277520 0 0 $X=2220238 $Y=2277118
X149 7451 4 6790 2 7478 NAND2X1 $T=2252580 2358160 0 0 $X=2252578 $Y=2357758
X150 7451 4 7477 2 7476 NAND2X1 $T=2260500 2358160 0 0 $X=2260498 $Y=2357758
X151 6790 4 7477 2 7479 NAND2X1 $T=2260500 2378320 1 0 $X=2260498 $Y=2372880
X152 7464 4 7512 2 7496 NAND2X1 $T=2270400 2297680 1 0 $X=2270398 $Y=2292240
X153 7643 4 7677 2 7675 NAND2X1 $T=2317920 2277520 1 0 $X=2317918 $Y=2272080
X154 7642 4 7651 2 7685 NAND2X1 $T=2319240 2307760 1 0 $X=2319238 $Y=2302320
X155 7685 4 7677 2 7706 NAND2X1 $T=2321220 2287600 1 180 $X=2319240 $Y=2287198
X156 7654 4 7818 2 7829 NAND2X1 $T=2356200 2307760 1 0 $X=2356198 $Y=2302320
X157 7847 4 7846 2 7859 NAND2X1 $T=2364120 2317840 1 180 $X=2362140 $Y=2317438
X158 7896 4 7946 2 8009 NAND2X1 $T=2408340 2267440 1 180 $X=2406360 $Y=2267038
X159 8083 4 8082 2 8101 NAND2X1 $T=2431440 2338000 1 180 $X=2429460 $Y=2337598
X160 8086 4 8083 2 8170 NAND2X1 $T=2440020 2338000 0 0 $X=2440018 $Y=2337598
X161 8199 4 8200 2 8219 NAND2X1 $T=2461800 2247280 0 0 $X=2461798 $Y=2246878
X162 8215 4 8186 2 8205 NAND2X1 $T=2466420 2287600 1 180 $X=2464440 $Y=2287198
X163 8287 4 8236 2 8309 NAND2X1 $T=2488200 2327920 0 180 $X=2486220 $Y=2322480
X164 8314 4 8283 2 8346 NAND2X1 $T=2496780 2287600 0 180 $X=2494800 $Y=2282160
X165 8309 4 8354 2 498 NAND2X1 $T=2509980 2247280 1 0 $X=2509978 $Y=2241840
X166 8463 4 8471 2 502 NAND2X1 $T=2528460 2257360 0 0 $X=2528458 $Y=2256958
X167 8505 4 8476 2 8490 NAND2X1 $T=2531760 2378320 0 180 $X=2529780 $Y=2372880
X168 8546 4 8549 2 8577 NAND2X1 $T=2544300 2317840 1 0 $X=2544298 $Y=2312400
X169 8475 4 8569 2 8525 NAND2X1 $T=2546940 2297680 0 0 $X=2546938 $Y=2297278
X170 8556 4 8611 2 8615 NAND2X1 $T=2557500 2338000 0 0 $X=2557498 $Y=2337598
X171 8614 4 8634 2 8599 NAND2X1 $T=2565420 2267440 0 0 $X=2565418 $Y=2267038
X172 8648 4 8666 2 8568 NAND2X1 $T=2573340 2287600 0 0 $X=2573338 $Y=2287198
X173 8574 4 8313 2 8729 NAND2X1 $T=2591820 2317840 1 0 $X=2591818 $Y=2312400
X174 2224 2 4 65 2242 NOR2X4 $T=911460 2257360 0 180 $X=906840 $Y=2251920
X175 2242 2 4 2330 2351 NOR2X4 $T=935880 2257360 1 0 $X=935878 $Y=2251920
X176 2332 2 4 66 2330 NOR2X4 $T=935880 2267440 0 0 $X=935878 $Y=2267038
X177 2807 2 4 1913 2808 NOR2X4 $T=1048740 2327920 0 0 $X=1048738 $Y=2327518
X178 2904 2 4 1815 2905 NOR2X4 $T=1079100 2358160 0 180 $X=1074480 $Y=2352720
X179 2906 2 4 1902 2908 NOR2X4 $T=1085040 2398480 0 180 $X=1080420 $Y=2393040
X180 3001 2 4 1609 2980 NOR2X4 $T=1104180 2338000 1 180 $X=1099560 $Y=2337598
X181 2905 2 4 2980 112 NOR2X4 $T=1100880 2368240 0 0 $X=1100878 $Y=2367838
X182 2908 2 4 2999 111 NOR2X4 $T=1105500 2398480 1 180 $X=1100880 $Y=2398078
X183 3640 2 4 2597 3712 NOR2X4 $T=1252680 2368240 0 0 $X=1252678 $Y=2367838
X184 2595 2 4 178 3917 NOR2X4 $T=1325280 2348080 0 180 $X=1320660 $Y=2342640
X185 288 2 4 2880 5217 NOR2X4 $T=1610400 2277520 1 0 $X=1610398 $Y=2272080
X186 351 2 4 3221 5857 NOR2X4 $T=1822260 2297680 1 180 $X=1817640 $Y=2297278
X187 382 2 4 3379 6314 NOR2X4 $T=1941060 2348080 1 180 $X=1936440 $Y=2347678
X188 7995 2 4 8072 8088 NOR2X4 $T=2429460 2277520 1 0 $X=2429458 $Y=2272080
X189 8201 2 4 8187 8217 NOR2X4 $T=2467740 2277520 0 180 $X=2463120 $Y=2272080
X190 1577 4 1558 1555 2 NAND2BX1 $T=711480 2307760 0 180 $X=708840 $Y=2302320
X191 1686 4 1684 1685 2 NAND2BX1 $T=749760 2327920 0 180 $X=747120 $Y=2322480
X192 1660 4 1669 1735 2 NAND2BX1 $T=749760 2338000 0 0 $X=749758 $Y=2337598
X193 50 4 49 1838 2 NAND2BX1 $T=789360 2267440 0 0 $X=789358 $Y=2267038
X194 1839 4 1687 1840 2 NAND2BX1 $T=793320 2358160 1 0 $X=793318 $Y=2352720
X195 51 4 52 1839 2 NAND2BX1 $T=796620 2348080 1 0 $X=796618 $Y=2342640
X196 2105 4 2088 2190 2 NAND2BX1 $T=875160 2348080 1 0 $X=875158 $Y=2342640
X197 2276 4 2309 2327 2 NAND2BX1 $T=927960 2348080 1 0 $X=927958 $Y=2342640
X198 2668 4 2652 2650 2 NAND2BX1 $T=1019040 2257360 1 180 $X=1016400 $Y=2256958
X199 2710 4 2713 2695 2 NAND2BX1 $T=1037520 2247280 1 180 $X=1034880 $Y=2246878
X200 2808 4 2769 2839 2 NAND2BX1 $T=1049400 2338000 0 0 $X=1049398 $Y=2337598
X201 2867 4 2842 2766 2 NAND2BX1 $T=1063260 2297680 0 180 $X=1060620 $Y=2292240
X202 3337 4 3311 3335 2 NAND2BX1 $T=1189320 2368240 1 0 $X=1189318 $Y=2362800
X203 149 4 3494 3478 2 NAND2BX1 $T=1218360 2267440 0 180 $X=1215720 $Y=2262000
X204 3483 4 3495 3545 2 NAND2BX1 $T=1222980 2358160 1 0 $X=1222978 $Y=2352720
X205 3299 4 3632 3633 2 NAND2BX1 $T=1246740 2297680 1 0 $X=1246738 $Y=2292240
X206 3596 4 3633 3624 2 NAND2BX1 $T=1246740 2297680 0 0 $X=1246738 $Y=2297278
X207 165 4 162 3682 2 NAND2BX1 $T=1257300 2237200 0 180 $X=1254660 $Y=2231760
X208 3667 4 3706 3754 2 NAND2BX1 $T=1261260 2338000 1 0 $X=1261258 $Y=2332560
X209 3683 4 3620 3804 2 NAND2BX1 $T=1266540 2358160 1 0 $X=1266538 $Y=2352720
X210 3712 4 3641 3831 2 NAND2BX1 $T=1279740 2368240 0 0 $X=1279738 $Y=2367838
X211 4028 4 4007 4008 2 NAND2BX1 $T=1343760 2388400 0 180 $X=1341120 $Y=2382960
X212 4102 4 4082 4100 2 NAND2BX1 $T=1370820 2378320 1 0 $X=1370818 $Y=2372880
X213 4145 4 4143 4140 2 NAND2BX1 $T=1374780 2327920 1 180 $X=1372140 $Y=2327518
X214 4230 4 4210 4182 2 NAND2BX1 $T=1394580 2257360 1 180 $X=1391940 $Y=2256958
X215 4231 4 4219 4215 2 NAND2BX1 $T=1397220 2287600 1 180 $X=1394580 $Y=2287198
X216 4654 4 4642 4641 2 NAND2BX1 $T=1503480 2247280 0 180 $X=1500840 $Y=2241840
X217 4719 4 4688 4644 2 NAND2BX1 $T=1519980 2388400 0 180 $X=1517340 $Y=2382960
X218 4779 4 4793 4802 2 NAND2BX1 $T=1543740 2277520 1 0 $X=1543738 $Y=2272080
X219 279 4 5095 5102 2 NAND2BX1 $T=1620960 2277520 0 0 $X=1620958 $Y=2277118
X220 5712 4 5707 5695 2 NAND2BX1 $T=1783320 2317840 1 180 $X=1780680 $Y=2317438
X221 5857 4 5927 5985 2 NAND2BX1 $T=1853940 2287600 1 0 $X=1853938 $Y=2282160
X222 6111 4 6108 6217 2 NAND2BX1 $T=1887600 2338000 1 0 $X=1887598 $Y=2332560
X223 6131 4 6133 6266 2 NAND2BX1 $T=1914000 2358160 0 0 $X=1913998 $Y=2357758
X224 6314 4 6322 6321 2 NAND2BX1 $T=1941060 2327920 0 180 $X=1938420 $Y=2322480
X225 6505 4 6534 399 2 NAND2BX1 $T=1993200 2317840 0 0 $X=1993198 $Y=2317438
X226 5244 4 6648 6634 2 NAND2BX1 $T=2023560 2297680 0 180 $X=2020920 $Y=2292240
X227 6802 4 6809 6857 2 NAND2BX1 $T=2070420 2307760 0 0 $X=2070418 $Y=2307358
X228 7035 4 7048 7066 2 NAND2BX1 $T=2143680 2247280 1 180 $X=2141040 $Y=2246878
X229 7039 4 7088 7114 2 NAND2BX1 $T=2162160 2257360 1 0 $X=2162158 $Y=2251920
X230 7448 4 7449 7396 2 NAND2BX1 $T=2253900 2257360 0 180 $X=2251260 $Y=2251920
X231 7482 4 7496 7508 2 NAND2BX1 $T=2270400 2267440 0 0 $X=2270398 $Y=2267038
X232 7828 4 7819 7817 2 NAND2BX1 $T=2358180 2287600 0 180 $X=2355540 $Y=2282160
X233 7862 4 7859 7861 2 NAND2BX1 $T=2370060 2297680 1 0 $X=2370058 $Y=2292240
X234 8187 4 8089 8200 2 NAND2BX1 $T=2460480 2267440 1 0 $X=2460478 $Y=2262000
X235 8201 4 8205 489 2 NAND2BX1 $T=2491500 2277520 1 0 $X=2491498 $Y=2272080
X236 8358 4 8346 490 2 NAND2BX1 $T=2502060 2267440 0 180 $X=2499420 $Y=2262000
X237 8461 4 8472 507 2 NAND2BX1 $T=2536380 2267440 0 0 $X=2536378 $Y=2267038
X238 8568 4 8569 8613 2 NAND2BX1 $T=2559480 2287600 0 0 $X=2559478 $Y=2287198
X239 1577 1572 4 1558 2 1593 OAI21X1 $T=724020 2307760 0 180 $X=720720 $Y=2302320
X240 1797 1643 4 1734 2 1799 OAI21X1 $T=780120 2317840 0 180 $X=776820 $Y=2312400
X241 1825 1687 4 1643 2 1818 OAI21X1 $T=788040 2317840 1 180 $X=784740 $Y=2317438
X242 2179 1899 4 2225 2 2329 OAI21X1 $T=915420 2348080 0 0 $X=915418 $Y=2347678
X243 3099 3023 4 3092 2 3094 OAI21X1 $T=1129920 2307760 0 180 $X=1126620 $Y=2302320
X244 3283 3337 4 3311 2 3328 OAI21X1 $T=1189980 2388400 0 180 $X=1186680 $Y=2382960
X245 3444 3483 4 3495 2 3498 OAI21X1 $T=1221660 2368240 0 180 $X=1218360 $Y=2362800
X246 3764 3712 4 3641 2 3720 OAI21X1 $T=1278420 2378320 1 0 $X=1278418 $Y=2372880
X247 4082 4028 4 4007 2 184 OAI21X1 $T=1355640 2388400 0 180 $X=1352340 $Y=2382960
X248 4221 4306 4 4309 2 207 OAI21X1 $T=1409100 2388400 0 0 $X=1409098 $Y=2387998
X249 267 4877 4 4880 2 4791 OAI21X1 $T=1560900 2237200 1 0 $X=1560898 $Y=2231760
X250 6361 374 4 6344 2 6356 OAI21X1 $T=1948320 2388400 1 180 $X=1945020 $Y=2387998
X251 7449 7482 4 7496 2 7498 OAI21X1 $T=2263800 2277520 0 0 $X=2263798 $Y=2277118
X252 8199 8201 4 8205 2 8249 OAI21X1 $T=2471700 2277520 1 0 $X=2471698 $Y=2272080
X253 8309 8358 4 8346 2 8357 OAI21X1 $T=2506680 2277520 0 180 $X=2503380 $Y=2272080
X254 1660 4 1668 1669 2 1723 OAI21XL $T=741840 2338000 1 0 $X=741838 $Y=2332560
X255 1669 4 1686 1684 2 1733 OAI21XL $T=748440 2317840 1 0 $X=748438 $Y=2312400
X256 1759 4 1687 1755 2 1757 OAI21XL $T=765600 2348080 1 180 $X=762960 $Y=2347678
X257 2088 4 2108 2107 2 2106 OAI21XL $T=873840 2338000 0 180 $X=871200 $Y=2332560
X258 2277 4 2309 2310 2 2240 OAI21XL $T=929280 2327920 1 180 $X=926640 $Y=2327518
X259 2276 4 2225 2309 2 2343 OAI21XL $T=927960 2358160 1 0 $X=927958 $Y=2352720
X260 2364 4 1899 2344 2 2425 OAI21XL $T=944460 2358160 1 0 $X=944458 $Y=2352720
X261 2413 4 1899 2442 2 2440 OAI21XL $T=962940 2358160 0 0 $X=962938 $Y=2357758
X262 2262 4 1899 2260 2 2519 OAI21XL $T=977460 2317840 0 0 $X=977458 $Y=2317438
X263 2520 4 1899 2500 2 2648 OAI21XL $T=989340 2307760 0 0 $X=989338 $Y=2307358
X264 2652 4 2710 2713 2 2696 OAI21XL $T=1029600 2257360 0 0 $X=1029598 $Y=2256958
X265 2716 4 2676 2672 2 2701 OAI21XL $T=1034880 2307760 0 180 $X=1032240 $Y=2302320
X266 2997 4 3091 3081 2 3098 OAI21XL $T=1126620 2267440 0 0 $X=1126618 $Y=2267038
X267 3152 4 3197 3204 2 3243 OAI21XL $T=1160940 2277520 1 0 $X=1160938 $Y=2272080
X268 3225 4 3023 3244 2 3254 OAI21XL $T=1162920 2317840 1 0 $X=1162918 $Y=2312400
X269 3219 4 3092 3294 2 3296 OAI21XL $T=1176120 2287600 1 0 $X=1176118 $Y=2282160
X270 3259 4 3309 3310 2 3274 OAI21XL $T=1181400 2297680 0 0 $X=1181398 $Y=2297278
X271 3270 4 3023 3275 2 3318 OAI21XL $T=1181400 2307760 0 0 $X=1181398 $Y=2307358
X272 3310 4 3334 3336 2 3255 OAI21XL $T=1188000 2277520 1 0 $X=1187998 $Y=2272080
X273 3326 4 140 3283 2 3355 OAI21XL $T=1195920 2408560 0 180 $X=1193280 $Y=2403120
X274 3426 4 140 3431 2 3472 OAI21XL $T=1203840 2398480 0 0 $X=1203838 $Y=2398078
X275 3477 4 3299 3471 2 3479 OAI21XL $T=1215720 2277520 1 0 $X=1215718 $Y=2272080
X276 3471 4 149 3494 2 3621 OAI21XL $T=1218360 2257360 1 0 $X=1218358 $Y=2251920
X277 3523 4 140 3499 2 3518 OAI21XL $T=1225620 2408560 0 180 $X=1222980 $Y=2403120
X278 3593 4 155 153 2 3625 OAI21XL $T=1238820 2237200 1 0 $X=1238818 $Y=2231760
X279 3665 4 3623 3666 2 3596 OAI21XL $T=1246740 2277520 0 180 $X=1244100 $Y=2272080
X280 157 4 140 3591 2 3690 OAI21XL $T=1246740 2408560 1 0 $X=1246738 $Y=2403120
X281 3668 4 3299 3623 2 3687 OAI21XL $T=1261260 2287600 1 180 $X=1258620 $Y=2287198
X282 3620 4 3667 3706 2 3675 OAI21XL $T=1259940 2348080 0 0 $X=1259938 $Y=2347678
X283 3753 4 3299 3718 2 3708 OAI21XL $T=1267860 2257360 0 180 $X=1265220 $Y=2251920
X284 3683 4 3724 3620 2 3749 OAI21XL $T=1267860 2368240 0 0 $X=1267858 $Y=2367838
X285 167 4 140 3745 2 3726 OAI21XL $T=1271820 2408560 1 180 $X=1269180 $Y=2408158
X286 165 4 3671 162 2 3763 OAI21XL $T=1273140 2237200 1 0 $X=1273138 $Y=2231760
X287 3742 4 3299 3810 2 3843 OAI21XL $T=1290300 2257360 0 0 $X=1290298 $Y=2256958
X288 3801 4 140 3827 2 3853 OAI21XL $T=1293600 2408560 1 0 $X=1293598 $Y=2403120
X289 3807 4 3299 3825 2 3882 OAI21XL $T=1295580 2257360 1 0 $X=1295578 $Y=2251920
X290 4145 4 4158 4143 2 4193 OAI21XL $T=1374780 2338000 1 0 $X=1374778 $Y=2332560
X291 4143 4 4213 4220 2 4216 OAI21XL $T=1394580 2327920 1 0 $X=1394578 $Y=2322480
X292 4234 4 4231 4219 2 4212 OAI21XL $T=1398540 2297680 1 180 $X=1395900 $Y=2297278
X293 4745 4 4737 4714 2 4734 OAI21XL $T=1531860 2327920 0 180 $X=1529220 $Y=2322480
X294 5062 4 290 5046 2 5100 OAI21XL $T=1615680 2388400 1 0 $X=1615678 $Y=2382960
X295 5046 4 5082 5098 2 293 OAI21XL $T=1627560 2378320 1 0 $X=1627558 $Y=2372880
X296 5137 4 290 5171 2 297 OAI21XL $T=1642080 2408560 0 0 $X=1642078 $Y=2408158
X297 310 4 5405 5404 2 5439 OAI21XL $T=1708740 2378320 0 0 $X=1708738 $Y=2377918
X298 295 4 321 5438 2 5470 OAI21XL $T=1716000 2247280 1 0 $X=1715998 $Y=2241840
X299 5464 4 5479 5481 2 327 OAI21XL $T=1725240 2398480 0 0 $X=1725238 $Y=2398078
X300 5481 4 5500 5504 2 5441 OAI21XL $T=1733160 2388400 0 0 $X=1733158 $Y=2387998
X301 5630 4 5348 5627 2 5629 OAI21XL $T=1764840 2358160 0 180 $X=1762200 $Y=2352720
X302 329 4 336 5650 2 5609 OAI21XL $T=1768800 2277520 1 0 $X=1768798 $Y=2272080
X303 5630 4 5348 5594 2 5717 OAI21XL $T=1779360 2358160 1 0 $X=1779358 $Y=2352720
X304 5754 4 5712 5707 2 5719 OAI21XL $T=1789260 2317840 0 180 $X=1786620 $Y=2312400
X305 5607 4 5348 5676 2 5817 OAI21XL $T=1805100 2358160 1 180 $X=1802460 $Y=2357758
X306 5676 4 5818 5724 2 5829 OAI21XL $T=1807740 2338000 1 180 $X=1805100 $Y=2337598
X307 5862 4 5348 5828 2 5889 OAI21XL $T=1819620 2338000 1 0 $X=1819618 $Y=2332560
X308 5888 4 5348 5890 2 5912 OAI21XL $T=1830180 2338000 0 0 $X=1830178 $Y=2337598
X309 6075 4 5993 6015 2 6120 OAI21XL $T=1884960 2398480 1 0 $X=1884958 $Y=2393040
X310 6108 4 6081 6028 2 6102 OAI21XL $T=1887600 2348080 1 180 $X=1884960 $Y=2347678
X311 6111 4 6138 6108 2 6218 OAI21XL $T=1892880 2358160 0 0 $X=1892878 $Y=2357758
X312 6131 4 6112 6133 2 6263 OAI21XL $T=1906080 2368240 1 0 $X=1906078 $Y=2362800
X313 6239 4 374 6192 2 6219 OAI21XL $T=1918620 2388400 1 180 $X=1915980 $Y=2387998
X314 6305 4 374 6286 2 6287 OAI21XL $T=1931820 2368240 1 180 $X=1929180 $Y=2367838
X315 6397 4 374 6398 2 6410 OAI21XL $T=1958220 2368240 0 0 $X=1958218 $Y=2367838
X316 7035 4 7053 7048 2 7113 OAI21XL $T=2147640 2247280 0 0 $X=2147638 $Y=2246878
X317 7048 4 7039 7088 2 7067 OAI21XL $T=2147640 2257360 1 0 $X=2147638 $Y=2251920
X318 8528 4 8525 8523 2 8519 OAI21XL $T=2541660 2287600 1 180 $X=2539020 $Y=2287198
X319 8568 4 8612 8528 2 8645 OAI21XL $T=2572680 2277520 1 180 $X=2570040 $Y=2277118
X320 8685 4 8612 8729 2 8681 OAI21XL $T=2581920 2277520 1 180 $X=2579280 $Y=2277118
X321 2293 2308 2328 4 2 XOR2X4 $T=924660 2297680 0 0 $X=924658 $Y=2297278
X322 2368 67 2455 4 2 XOR2X4 $T=945780 2297680 0 0 $X=945778 $Y=2297278
X323 2482 83 2504 4 2 XOR2X4 $T=975480 2287600 0 0 $X=975478 $Y=2287198
X324 87 2522 2595 4 2 XOR2X4 $T=989340 2267440 0 0 $X=989338 $Y=2267038
X325 2669 2664 2735 4 2 XOR2X4 $T=1020360 2398480 0 0 $X=1020358 $Y=2398078
X326 2723 2738 95 4 2 XOR2X4 $T=1034880 2408560 0 0 $X=1034878 $Y=2408158
X327 2839 2847 2880 4 2 XOR2X4 $T=1060620 2338000 0 0 $X=1060618 $Y=2337598
X328 3046 3074 3159 4 2 XOR2X4 $T=1115400 2358160 0 0 $X=1115398 $Y=2357758
X329 3077 3106 3256 4 2 XOR2X4 $T=1123980 2348080 0 0 $X=1123978 $Y=2347678
X330 3100 3203 3221 4 2 XOR2X4 $T=1147740 2398480 0 0 $X=1147738 $Y=2398078
X331 3335 3362 3379 4 2 XOR2X4 $T=1188000 2368240 0 0 $X=1187998 $Y=2367838
X332 3545 3473 3669 4 2 XOR2X4 $T=1228260 2358160 1 0 $X=1228258 $Y=2352720
X333 3546 3566 3670 4 2 XOR2X4 $T=1228260 2388400 1 0 $X=1228258 $Y=2382960
X334 3754 3782 169 4 2 XOR2X4 $T=1276440 2338000 1 0 $X=1276438 $Y=2332560
X335 3831 174 3896 4 2 XOR2X4 $T=1296240 2368240 0 0 $X=1296238 $Y=2367838
X336 3804 3899 190 4 2 XOR2X4 $T=1302840 2358160 1 0 $X=1302838 $Y=2352720
X337 3958 3976 183 4 2 XOR2X4 $T=1326600 2307760 1 0 $X=1326598 $Y=2302320
X338 4399 4420 225 4 2 XOR2X4 $T=1446720 2358160 0 0 $X=1446718 $Y=2357758
X339 4533 4472 239 4 2 XOR2X4 $T=1475760 2368240 0 0 $X=1475758 $Y=2367838
X340 277 5230 5244 4 2 XOR2X4 $T=1650660 2277520 1 0 $X=1650658 $Y=2272080
X341 6006 6023 361 4 2 XOR2X4 $T=1858560 2247280 1 0 $X=1858558 $Y=2241840
X342 6057 6077 364 4 2 XOR2X4 $T=1871760 2267440 1 0 $X=1871758 $Y=2262000
X343 6237 6265 378 4 2 XOR2X4 $T=1918620 2267440 1 0 $X=1918618 $Y=2262000
X344 6285 6262 381 4 2 XOR2X4 $T=1927860 2277520 1 0 $X=1927858 $Y=2272080
X345 6486 6465 388 4 2 XOR2X4 $T=1980660 2287600 1 180 $X=1969440 $Y=2287198
X346 6508 6633 407 4 2 XOR2X4 $T=2011020 2237200 1 0 $X=2011018 $Y=2231760
X347 338 5897 6731 4 2 XOR2X4 $T=2011680 2378320 1 0 $X=2011678 $Y=2372880
X348 1622 4 2 1625 INVX1 $T=729960 2317840 0 0 $X=729958 $Y=2317438
X349 1593 4 2 1668 INVX1 $T=737220 2327920 1 0 $X=737218 $Y=2322480
X350 1643 4 2 1756 INVX1 $T=767580 2327920 0 180 $X=766260 $Y=2322480
X351 1783 4 2 1871 INVX1 $T=787380 2297680 1 0 $X=787378 $Y=2292240
X352 1839 4 2 1850 INVX1 $T=799260 2348080 1 0 $X=799258 $Y=2342640
X353 1796 4 2 1847 INVX1 $T=799920 2277520 0 0 $X=799918 $Y=2277118
X354 2145 4 2 2151 INVX1 $T=886380 2338000 1 0 $X=886378 $Y=2332560
X355 2174 4 2 2148 INVX1 $T=890340 2338000 1 180 $X=889020 $Y=2337598
X356 2106 4 2 2167 INVX1 $T=892980 2338000 0 180 $X=891660 $Y=2332560
X357 2294 4 2 2313 INVX1 $T=932580 2287600 0 180 $X=931260 $Y=2282160
X358 2330 4 2 2318 INVX1 $T=937200 2277520 1 180 $X=935880 $Y=2277118
X359 2380 4 2 2346 INVX1 $T=945780 2348080 0 180 $X=944460 $Y=2342640
X360 2355 4 2 2413 INVX1 $T=953700 2358160 0 0 $X=953698 $Y=2357758
X361 2438 4 2 2354 INVX1 $T=955680 2338000 0 180 $X=954360 $Y=2332560
X362 68 4 2 2454 INVX1 $T=955680 2257360 0 0 $X=955678 $Y=2256958
X363 2343 4 2 2442 INVX1 $T=962280 2358160 1 0 $X=962278 $Y=2352720
X364 78 4 2 2488 INVX1 $T=966240 2267440 1 0 $X=966238 $Y=2262000
X365 2598 4 2 2599 INVX1 $T=1009140 2388400 1 0 $X=1009138 $Y=2382960
X366 2633 4 2 2693 INVX1 $T=1022340 2398480 1 0 $X=1022338 $Y=2393040
X367 2731 4 2 2734 INVX1 $T=1038180 2378320 1 0 $X=1038178 $Y=2372880
X368 2740 4 2 2751 INVX1 $T=1052700 2398480 0 180 $X=1051380 $Y=2393040
X369 2867 4 2 2878 INVX1 $T=1069860 2297680 1 0 $X=1069858 $Y=2292240
X370 2999 4 2 3107 INVX1 $T=1124640 2408560 0 0 $X=1124638 $Y=2408158
X371 3092 4 2 3198 INVX1 $T=1150380 2297680 0 0 $X=1150378 $Y=2297278
X372 3099 4 2 3224 INVX1 $T=1158300 2297680 0 0 $X=1158298 $Y=2297278
X373 2616 4 2 134 INVX1 $T=1182720 2408560 0 0 $X=1182718 $Y=2408158
X374 3326 4 2 3317 INVX1 $T=1186020 2398480 0 180 $X=1184700 $Y=2393040
X375 3450 4 2 3432 INVX1 $T=1207140 2287600 1 180 $X=1205820 $Y=2287198
X376 3444 4 2 3430 INVX1 $T=1212420 2388400 0 180 $X=1211100 $Y=2382960
X377 3328 4 2 3499 INVX1 $T=1216380 2398480 1 0 $X=1216378 $Y=2393040
X378 3299 4 2 3475 INVX1 $T=1219680 2297680 1 0 $X=1219678 $Y=2292240
X379 3517 4 2 3425 INVX1 $T=1222980 2378320 1 180 $X=1221660 $Y=2377918
X380 3333 4 2 3523 INVX1 $T=1223640 2398480 0 0 $X=1223638 $Y=2398078
X381 3621 4 2 3623 INVX1 $T=1244760 2257360 1 0 $X=1244758 $Y=2251920
X382 3665 4 2 3672 INVX1 $T=1252680 2267440 0 0 $X=1252678 $Y=2267038
X383 161 4 2 163 INVX1 $T=1255320 2408560 0 0 $X=1255318 $Y=2408158
X384 3623 4 2 3691 INVX1 $T=1257960 2257360 1 0 $X=1257958 $Y=2251920
X385 3591 4 2 166 INVX1 $T=1267860 2398480 1 0 $X=1267858 $Y=2393040
X386 3671 4 2 3747 INVX1 $T=1268520 2237200 1 0 $X=1268518 $Y=2231760
X387 157 4 2 3752 INVX1 $T=1268520 2408560 1 0 $X=1268518 $Y=2403120
X388 3720 4 2 3724 INVX1 $T=1269840 2378320 0 180 $X=1268520 $Y=2372880
X389 3741 4 2 3751 INVX1 $T=1271160 2247280 1 0 $X=1271158 $Y=2241840
X390 3526 4 2 3668 INVX1 $T=1272480 2287600 0 180 $X=1271160 $Y=2282160
X391 3695 4 2 3725 INVX1 $T=1272480 2388400 1 180 $X=1271160 $Y=2387998
X392 3766 4 2 3788 INVX1 $T=1284360 2388400 1 0 $X=1284358 $Y=2382960
X393 3880 4 2 3883 INVX1 $T=1303500 2297680 1 0 $X=1303498 $Y=2292240
X394 3881 4 2 3929 INVX1 $T=1311420 2287600 0 0 $X=1311418 $Y=2287198
X395 3914 4 2 3961 INVX1 $T=1315380 2317840 0 0 $X=1315378 $Y=2317438
X396 3898 4 2 3916 INVX1 $T=1319340 2247280 1 180 $X=1318020 $Y=2246878
X397 3917 4 2 3993 INVX1 $T=1339140 2338000 0 0 $X=1339138 $Y=2337598
X398 4082 4 2 4070 INVX1 $T=1355640 2378320 0 180 $X=1354320 $Y=2372880
X399 4067 4 2 4119 INVX1 $T=1355640 2327920 1 0 $X=1355638 $Y=2322480
X400 4085 4 2 4118 INVX1 $T=1370160 2297680 1 0 $X=1370158 $Y=2292240
X401 4013 4 2 4137 INVX1 $T=1378080 2307760 0 0 $X=1378078 $Y=2307358
X402 4212 4 2 4158 INVX1 $T=1389960 2338000 1 180 $X=1388640 $Y=2337598
X403 205 4 2 4314 INVX1 $T=1407120 2297680 0 0 $X=1407118 $Y=2297278
X404 4279 4 2 4276 INVX1 $T=1409760 2368240 0 0 $X=1409758 $Y=2367838
X405 201 4 2 206 INVX1 $T=1410420 2237200 0 0 $X=1410418 $Y=2236798
X406 4295 4 2 4229 INVX1 $T=1417680 2247280 1 180 $X=1416360 $Y=2246878
X407 4330 4 2 4343 INVX1 $T=1420320 2368240 1 0 $X=1420318 $Y=2362800
X408 4538 4 2 4491 INVX1 $T=1479720 2378320 1 0 $X=1479718 $Y=2372880
X409 4733 4 2 4660 INVX1 $T=1528560 2378320 0 180 $X=1527240 $Y=2372880
X410 4755 4 2 4705 INVX1 $T=1529880 2287600 1 180 $X=1528560 $Y=2287198
X411 4756 4 2 4766 INVX1 $T=1537800 2317840 1 0 $X=1537798 $Y=2312400
X412 4852 4 2 4768 INVX1 $T=1549680 2257360 1 180 $X=1548360 $Y=2256958
X413 5033 4 2 5031 INVX1 $T=1611060 2237200 0 0 $X=1611058 $Y=2236798
X414 281 4 2 5095 INVX1 $T=1622280 2237200 1 0 $X=1622278 $Y=2231760
X415 5231 4 2 5247 INVX1 $T=1663200 2267440 0 0 $X=1663198 $Y=2267038
X416 5260 4 2 5259 INVX1 $T=1669800 2378320 0 180 $X=1668480 $Y=2372880
X417 301 4 2 5283 INVX1 $T=1673760 2408560 0 0 $X=1673758 $Y=2408158
X418 5328 4 2 5294 INVX1 $T=1688280 2398480 0 180 $X=1686960 $Y=2393040
X419 316 4 2 5345 INVX1 $T=1702140 2257360 1 0 $X=1702138 $Y=2251920
X420 5395 4 2 5443 INVX1 $T=1716000 2398480 1 0 $X=1715998 $Y=2393040
X421 5439 4 2 5479 INVX1 $T=1720620 2398480 0 0 $X=1720618 $Y=2398078
X422 271 4 2 5517 INVX1 $T=1736460 2287600 0 0 $X=1736458 $Y=2287198
X423 260 4 2 333 INVX1 $T=1749660 2247280 0 180 $X=1748340 $Y=2241840
X424 5609 4 2 5647 INVX1 $T=1760220 2267440 1 0 $X=1760218 $Y=2262000
X425 314 4 2 5150 INVX1 $T=1760220 2297680 0 0 $X=1760218 $Y=2297278
X426 5651 4 2 5671 INVX1 $T=1770120 2388400 0 0 $X=1770118 $Y=2387998
X427 5655 4 2 5818 INVX1 $T=1797180 2338000 0 0 $X=1797178 $Y=2337598
X428 5737 4 2 5847 INVX1 $T=1804440 2317840 0 0 $X=1804438 $Y=2317438
X429 338 4 2 345 INVX1 $T=1816320 2388400 1 180 $X=1815000 $Y=2387998
X430 348 4 2 320 INVX1 $T=1818960 2247280 0 0 $X=1818958 $Y=2246878
X431 5858 4 2 5888 INVX1 $T=1820940 2338000 0 0 $X=1820938 $Y=2337598
X432 5829 4 2 5890 INVX1 $T=1825560 2338000 0 0 $X=1825558 $Y=2337598
X433 5924 4 2 5891 INVX1 $T=1832160 2388400 0 180 $X=1830840 $Y=2382960
X434 321 4 2 349 INVX1 $T=1861860 2408560 1 0 $X=1861858 $Y=2403120
X435 6061 4 2 6078 INVX1 $T=1875060 2297680 0 0 $X=1875058 $Y=2297278
X436 6120 4 2 6138 INVX1 $T=1894860 2368240 0 180 $X=1893540 $Y=2362800
X437 6189 4 2 6151 INVX1 $T=1900140 2287600 0 180 $X=1898820 $Y=2282160
X438 6140 4 2 6222 INVX1 $T=1906080 2408560 1 0 $X=1906078 $Y=2403120
X439 6075 4 2 6252 INVX1 $T=1914660 2408560 0 0 $X=1914658 $Y=2408158
X440 6234 4 2 6254 INVX1 $T=1917300 2317840 1 0 $X=1917298 $Y=2312400
X441 6259 4 2 6237 INVX1 $T=1923900 2267440 1 180 $X=1922580 $Y=2267038
X442 6112 4 2 6277 INVX1 $T=1925220 2358160 0 0 $X=1925218 $Y=2357758
X443 6202 4 2 6269 INVX1 $T=1933800 2368240 0 0 $X=1933798 $Y=2367838
X444 370 4 2 6344 INVX1 $T=1941720 2388400 1 180 $X=1940400 $Y=2387998
X445 375 4 2 6361 INVX1 $T=1947000 2398480 0 0 $X=1946998 $Y=2398078
X446 374 4 2 376 INVX1 $T=1952280 2408560 1 0 $X=1952278 $Y=2403120
X447 6474 4 2 6467 INVX1 $T=1976040 2327920 1 180 $X=1974720 $Y=2327518
X448 6449 4 2 6500 INVX1 $T=1980000 2247280 1 0 $X=1979998 $Y=2241840
X449 6501 4 2 396 INVX1 $T=1985940 2257360 0 0 $X=1985938 $Y=2256958
X450 6634 4 2 6650 INVX1 $T=2018940 2287600 0 0 $X=2018938 $Y=2287198
X451 5244 4 2 6662 INVX1 $T=2021580 2327920 1 0 $X=2021578 $Y=2322480
X452 6678 4 2 6693 INVX1 $T=2032140 2398480 0 0 $X=2032138 $Y=2398078
X453 5266 4 2 6691 INVX1 $T=2044680 2327920 1 0 $X=2044678 $Y=2322480
X454 5106 4 2 6709 INVX1 $T=2046000 2317840 1 180 $X=2044680 $Y=2317438
X455 6805 4 2 6825 INVX1 $T=2071080 2327920 0 0 $X=2071078 $Y=2327518
X456 6787 4 2 6809 INVX1 $T=2072400 2297680 1 180 $X=2071080 $Y=2297278
X457 5988 4 2 6868 INVX1 $T=2087580 2398480 0 180 $X=2086260 $Y=2393040
X458 6857 4 2 6863 INVX1 $T=2086920 2297680 0 0 $X=2086918 $Y=2297278
X459 6858 4 2 6886 INVX1 $T=2086920 2317840 0 0 $X=2086918 $Y=2317438
X460 6854 4 2 6877 INVX1 $T=2092200 2297680 0 0 $X=2092198 $Y=2297278
X461 6958 4 2 6961 INVX1 $T=2105400 2358160 0 0 $X=2105398 $Y=2357758
X462 6962 4 2 427 INVX1 $T=2112660 2408560 1 0 $X=2112658 $Y=2403120
X463 431 4 2 6980 INVX1 $T=2119920 2257360 1 180 $X=2118600 $Y=2256958
X464 7166 4 2 7229 INVX1 $T=2173380 2267440 1 0 $X=2173378 $Y=2262000
X465 447 4 2 445 INVX1 $T=2183280 2408560 1 180 $X=2181960 $Y=2408158
X466 7303 4 2 7304 INVX1 $T=2216280 2267440 1 180 $X=2214960 $Y=2267038
X467 7685 4 2 7674 INVX1 $T=2321220 2297680 1 180 $X=2319900 $Y=2297278
X468 470 4 2 468 INVX1 $T=2397120 2237200 0 180 $X=2395800 $Y=2231760
X469 8039 4 2 8099 INVX1 $T=2442660 2247280 1 0 $X=2442658 $Y=2241840
X470 8187 4 2 8176 INVX1 $T=2454540 2257360 0 180 $X=2453220 $Y=2251920
X471 8309 4 2 8345 INVX1 $T=2497440 2247280 1 0 $X=2497438 $Y=2241840
X472 8353 4 2 8354 INVX1 $T=2502720 2247280 0 0 $X=2502718 $Y=2246878
X473 8463 4 2 8609 INVX1 $T=2552880 2267440 0 0 $X=2552878 $Y=2267038
X474 8357 4 2 8612 INVX1 $T=2552880 2277520 0 0 $X=2552878 $Y=2277118
X475 8577 4 2 8516 INVX1 $T=2552880 2307760 1 0 $X=2552878 $Y=2302320
X476 8528 4 2 8618 INVX1 $T=2566740 2297680 1 180 $X=2565420 $Y=2297278
X477 8615 4 2 8647 INVX1 $T=2578620 2307760 1 0 $X=2578618 $Y=2302320
X478 8685 4 2 8666 INVX1 $T=2582580 2287600 1 180 $X=2581260 $Y=2287198
X479 8729 4 2 8649 INVX1 $T=2593140 2297680 1 180 $X=2591820 $Y=2297278
X480 74 73 2 69 72 4 AOI21X2 $T=955020 2237200 0 180 $X=950400 $Y=2231760
X481 2696 2697 2 2701 2737 4 AOI21X2 $T=1027620 2287600 0 0 $X=1027618 $Y=2287198
X482 2616 2845 2 2840 2847 4 AOI21X2 $T=1065900 2378320 0 180 $X=1061280 $Y=2372880
X483 2616 3059 2 3039 3074 4 AOI21X2 $T=1117380 2368240 1 0 $X=1117378 $Y=2362800
X484 2616 124 2 3035 3203 4 AOI21X2 $T=1152360 2408560 0 180 $X=1147740 $Y=2403120
X485 132 3363 2 3355 3362 4 AOI21X2 $T=1196580 2408560 1 180 $X=1191960 $Y=2408158
X486 132 3446 2 3472 3473 4 AOI21X2 $T=1215060 2408560 0 180 $X=1210440 $Y=2403120
X487 3516 3328 2 3498 3591 4 AOI21X2 $T=1221660 2398480 1 0 $X=1221658 $Y=2393040
X488 164 132 2 3690 3709 4 AOI21X2 $T=1264560 2408560 0 180 $X=1259940 $Y=2403120
X489 168 132 2 3726 3782 4 AOI21X2 $T=1283700 2408560 1 180 $X=1279080 $Y=2408158
X490 177 3883 2 3929 3928 4 AOI21X2 $T=1315380 2277520 1 0 $X=1315378 $Y=2272080
X491 4067 4086 2 4118 4160 4 AOI21X2 $T=1362240 2287600 0 0 $X=1362238 $Y=2287198
X492 4118 4066 2 4137 4124 4 AOI21X2 $T=1368180 2307760 1 0 $X=1368178 $Y=2302320
X493 4755 4754 2 4734 4746 4 AOI21X2 $T=1537140 2327920 1 180 $X=1532520 $Y=2327518
X494 4791 4776 2 4768 4764 4 AOI21X2 $T=1541760 2257360 1 180 $X=1537140 $Y=2256958
X495 5329 5264 2 5346 5348 4 AOI21X2 $T=1692240 2388400 1 0 $X=1692238 $Y=2382960
X496 6509 6444 2 6467 6472 4 AOI21X2 $T=1976700 2327920 0 180 $X=1972080 $Y=2322480
X497 392 6473 2 6509 6465 4 AOI21X2 $T=1983300 2297680 1 0 $X=1983298 $Y=2292240
X498 6877 6864 2 6886 6897 4 AOI21X2 $T=2096820 2327920 0 180 $X=2092200 $Y=2322480
X499 7009 7054 2 7067 7086 4 AOI21X2 $T=2139060 2257360 1 0 $X=2139058 $Y=2251920
X500 7677 7671 2 7674 7689 4 AOI21X2 $T=2322540 2287600 0 180 $X=2317920 $Y=2282160
X501 478 8099 2 8103 479 4 AOI21X2 $T=2435400 2237200 1 0 $X=2435398 $Y=2231760
X502 478 8122 2 8089 482 4 AOI21X2 $T=2457840 2257360 1 0 $X=2457838 $Y=2251920
X503 8216 478 2 8219 485 4 AOI21X2 $T=2470380 2237200 1 180 $X=2465760 $Y=2236798
X504 8354 493 2 8345 494 4 AOI21X2 $T=2503380 2237200 0 180 $X=2498760 $Y=2231760
X505 2 1559 1543 1577 4 NOR2X1 $T=714780 2297680 0 0 $X=714778 $Y=2297278
X506 2 1610 32 1622 4 NOR2X1 $T=720720 2297680 1 0 $X=720718 $Y=2292240
X507 2 1577 1622 1638 4 NOR2X1 $T=730620 2307760 1 0 $X=730618 $Y=2302320
X508 2 1574 1657 1660 4 NOR2X1 $T=740520 2297680 0 0 $X=740518 $Y=2297278
X509 2 1686 1660 1737 4 NOR2X1 $T=749760 2307760 0 180 $X=747780 $Y=2302320
X510 2 1736 1673 1686 4 NOR2X1 $T=762960 2297680 0 180 $X=760980 $Y=2292240
X511 2 50 51 1783 4 NOR2X1 $T=787380 2277520 0 0 $X=787378 $Y=2277118
X512 2 1797 1825 1876 4 NOR2X1 $T=787380 2317840 1 0 $X=787378 $Y=2312400
X513 2 2076 1738 2105 4 NOR2X1 $T=865260 2327920 1 0 $X=865258 $Y=2322480
X514 2 2059 2089 2108 4 NOR2X1 $T=874500 2307760 1 0 $X=874498 $Y=2302320
X515 2 2108 2105 2174 4 NOR2X1 $T=877140 2327920 1 0 $X=877138 $Y=2322480
X516 2 2277 2276 2189 4 NOR2X1 $T=919380 2327920 1 180 $X=917400 $Y=2327518
X517 2 2276 2179 2355 4 NOR2X1 $T=919380 2358160 1 180 $X=917400 $Y=2357758
X518 2 2296 2172 2276 4 NOR2X1 $T=920700 2317840 1 180 $X=918720 $Y=2317438
X519 2 93 92 2668 4 NOR2X1 $T=1024320 2237200 0 180 $X=1022340 $Y=2231760
X520 2 2676 2689 2697 4 NOR2X1 $T=1025640 2297680 0 0 $X=1025638 $Y=2297278
X521 2 2674 2690 2689 4 NOR2X1 $T=1028280 2327920 0 180 $X=1026300 $Y=2322480
X522 2 2668 2710 2699 4 NOR2X1 $T=1037520 2257360 0 0 $X=1037518 $Y=2256958
X523 2 96 2765 2710 4 NOR2X1 $T=1047420 2257360 0 180 $X=1045440 $Y=2251920
X524 2 2866 2809 2676 4 NOR2X1 $T=1052040 2277520 0 180 $X=1050060 $Y=2272080
X525 2 2919 2867 2974 4 NOR2X1 $T=1084380 2297680 1 0 $X=1084378 $Y=2292240
X526 2 103 2937 2919 4 NOR2X1 $T=1087680 2267440 0 180 $X=1085700 $Y=2262000
X527 2 2918 2922 2867 4 NOR2X1 $T=1089660 2277520 0 0 $X=1089658 $Y=2277118
X528 2 2980 3024 3059 4 NOR2X1 $T=1111440 2378320 0 180 $X=1109460 $Y=2372880
X529 2 114 115 3003 4 NOR2X1 $T=1111440 2267440 0 0 $X=1111438 $Y=2267038
X530 2 2999 99 3101 4 NOR2X1 $T=1123980 2408560 1 0 $X=1123978 $Y=2403120
X531 2 3091 3003 3082 4 NOR2X1 $T=1125960 2277520 1 180 $X=1123980 $Y=2277118
X532 2 119 3083 3091 4 NOR2X1 $T=1135200 2257360 0 180 $X=1133220 $Y=2251920
X533 2 3126 120 3146 4 NOR2X1 $T=1137180 2267440 1 0 $X=1137178 $Y=2262000
X534 2 3197 3146 3218 4 NOR2X1 $T=1149060 2277520 0 0 $X=1149058 $Y=2277118
X535 2 3219 3099 3292 4 NOR2X1 $T=1160940 2287600 0 0 $X=1160938 $Y=2287198
X536 2 128 127 3197 4 NOR2X1 $T=1173480 2247280 0 180 $X=1171500 $Y=2241840
X537 2 133 130 3259 4 NOR2X1 $T=1180740 2257360 0 180 $X=1178760 $Y=2251920
X538 2 3334 3259 3220 4 NOR2X1 $T=1184040 2277520 1 180 $X=1182060 $Y=2277118
X539 2 136 137 3334 4 NOR2X1 $T=1191300 2247280 1 180 $X=1189320 $Y=2246878
X540 2 3326 143 3363 4 NOR2X1 $T=1202520 2408560 0 0 $X=1202518 $Y=2408158
X541 2 3426 143 3446 4 NOR2X1 $T=1205160 2408560 1 0 $X=1205158 $Y=2403120
X542 2 144 145 3477 4 NOR2X1 $T=1210440 2257360 1 0 $X=1210438 $Y=2251920
X543 2 149 3477 3526 4 NOR2X1 $T=1223640 2257360 1 0 $X=1223638 $Y=2251920
X544 2 154 152 3611 4 NOR2X1 $T=1239480 2267440 1 0 $X=1239478 $Y=2262000
X545 2 3523 143 3592 4 NOR2X1 $T=1239480 2408560 1 0 $X=1239478 $Y=2403120
X546 2 155 3611 3627 4 NOR2X1 $T=1244760 2247280 1 0 $X=1244758 $Y=2241840
X547 2 159 158 3665 4 NOR2X1 $T=1247400 2257360 0 0 $X=1247398 $Y=2256958
X548 2 3665 3668 3632 4 NOR2X1 $T=1254660 2287600 0 180 $X=1252680 $Y=2282160
X549 2 3667 3683 3684 4 NOR2X1 $T=1255320 2358160 1 0 $X=1255318 $Y=2352720
X550 2 3683 3725 3728 4 NOR2X1 $T=1267860 2388400 0 0 $X=1267858 $Y=2387998
X551 2 3794 2648 3880 4 NOR2X1 $T=1293600 2297680 1 0 $X=1293598 $Y=2292240
X552 2 3801 143 3886 4 NOR2X1 $T=1300860 2408560 1 0 $X=1300858 $Y=2403120
X553 2 176 2504 3914 4 NOR2X1 $T=1309440 2317840 1 180 $X=1307460 $Y=2317438
X554 2 4028 4102 189 4 NOR2X1 $T=1362900 2388400 1 0 $X=1362898 $Y=2382960
X555 2 4183 4180 4102 4 NOR2X1 $T=1385340 2378320 0 180 $X=1383360 $Y=2372880
X556 2 4213 4145 4214 4 NOR2X1 $T=1393260 2327920 1 180 $X=1391280 $Y=2327518
X557 2 201 196 4231 4 NOR2X1 $T=1398540 2277520 0 180 $X=1396560 $Y=2272080
X558 2 209 4314 4213 4 NOR2X1 $T=1417020 2327920 0 180 $X=1415040 $Y=2322480
X559 2 4382 197 4295 4 NOR2X1 $T=1435500 2247280 1 180 $X=1433520 $Y=2246878
X560 2 4464 4462 226 4 NOR2X1 $T=1457280 2408560 0 0 $X=1457278 $Y=2408158
X561 2 212 4645 4654 4 NOR2X1 $T=1504800 2267440 0 0 $X=1504798 $Y=2267038
X562 2 4756 4705 4711 4 NOR2X1 $T=1527900 2297680 1 180 $X=1525920 $Y=2297278
X563 2 4756 4737 4754 4 NOR2X1 $T=1537140 2327920 1 0 $X=1537138 $Y=2322480
X564 2 4777 4781 4733 4 NOR2X1 $T=1542420 2368240 0 180 $X=1540440 $Y=2362800
X565 2 4794 4789 4756 4 NOR2X1 $T=1543740 2297680 1 180 $X=1541760 $Y=2297278
X566 2 4882 4824 4779 4 NOR2X1 $T=1559580 2277520 1 180 $X=1557600 $Y=2277118
X567 2 4952 4901 4877 4 NOR2X1 $T=1573440 2237200 0 180 $X=1571460 $Y=2231760
X568 2 4708 5048 5062 4 NOR2X1 $T=1609080 2358160 1 0 $X=1609078 $Y=2352720
X569 2 5082 5062 5069 4 NOR2X1 $T=1617660 2378320 0 180 $X=1615680 $Y=2372880
X570 2 5068 5096 5082 4 NOR2X1 $T=1622940 2348080 1 180 $X=1620960 $Y=2347678
X571 2 5313 5312 308 4 NOR2X1 $T=1686960 2368240 0 180 $X=1684980 $Y=2362800
X572 2 5328 306 5329 4 NOR2X1 $T=1696200 2398480 1 180 $X=1694220 $Y=2398078
X573 2 5405 308 5395 4 NOR2X1 $T=1706100 2388400 1 180 $X=1704120 $Y=2387998
X574 2 5406 5323 5405 4 NOR2X1 $T=1709400 2348080 1 180 $X=1707420 $Y=2347678
X575 2 5500 5464 5426 4 NOR2X1 $T=1722600 2398480 0 180 $X=1720620 $Y=2393040
X576 2 5464 5443 325 4 NOR2X1 $T=1725240 2408560 1 180 $X=1723260 $Y=2408158
X577 2 5524 5422 5464 4 NOR2X1 $T=1735800 2398480 1 180 $X=1733820 $Y=2398078
X578 2 5519 5523 5500 4 NOR2X1 $T=1741740 2368240 0 0 $X=1741738 $Y=2367838
X579 2 5601 5546 5607 4 NOR2X1 $T=1756260 2338000 0 0 $X=1756258 $Y=2337598
X580 2 5712 5737 5713 4 NOR2X1 $T=1788600 2317840 0 0 $X=1788598 $Y=2317438
X581 2 5818 5607 5858 4 NOR2X1 $T=1816980 2338000 0 0 $X=1816978 $Y=2337598
X582 2 5833 5931 5993 4 NOR2X1 $T=1851300 2388400 0 0 $X=1851298 $Y=2387998
X583 2 6045 5910 6111 4 NOR2X1 $T=1869780 2338000 1 0 $X=1869778 $Y=2332560
X584 2 6034 5863 6081 4 NOR2X1 $T=1871760 2348080 0 0 $X=1871758 $Y=2347678
X585 2 5986 5830 6140 4 NOR2X1 $T=1877700 2398480 0 0 $X=1877698 $Y=2398078
X586 2 365 5645 6131 4 NOR2X1 $T=1888260 2368240 0 0 $X=1888258 $Y=2367838
X587 2 6081 6111 6116 4 NOR2X1 $T=1892880 2348080 0 0 $X=1892878 $Y=2347678
X588 2 5993 6140 6142 4 NOR2X1 $T=1894200 2388400 0 0 $X=1894198 $Y=2387998
X589 2 6131 6202 6267 4 NOR2X1 $T=1916640 2368240 0 0 $X=1916638 $Y=2367838
X590 2 6304 4065 6442 4 NOR2X1 $T=1956900 2267440 0 0 $X=1956898 $Y=2267038
X591 2 6500 6431 6508 4 NOR2X1 $T=1983300 2237200 0 0 $X=1983298 $Y=2236798
X592 2 6694 6710 6713 4 NOR2X1 $T=2044680 2277520 0 0 $X=2044678 $Y=2277118
X593 2 6947 6980 6992 4 NOR2X1 $T=2112660 2277520 0 180 $X=2110680 $Y=2272080
X594 2 430 6994 7035 4 NOR2X1 $T=2117940 2247280 0 0 $X=2117938 $Y=2246878
X595 2 7035 7039 7054 4 NOR2X1 $T=2133120 2257360 1 0 $X=2133118 $Y=2251920
X596 2 7071 7138 441 4 NOR2X1 $T=2168760 2408560 0 0 $X=2168758 $Y=2408158
X597 2 7448 7482 7484 4 NOR2X1 $T=2262480 2267440 0 0 $X=2262478 $Y=2267038
X598 2 7896 7946 8039 4 NOR2X1 $T=2406360 2267440 1 0 $X=2406358 $Y=2262000
X599 2 8287 8236 8353 4 NOR2X1 $T=2492160 2327920 1 0 $X=2492158 $Y=2322480
X600 2 8314 8283 8358 4 NOR2X1 $T=2499420 2287600 1 0 $X=2499418 $Y=2282160
X601 2 8358 8353 8463 4 NOR2X1 $T=2510640 2267440 1 0 $X=2510638 $Y=2262000
X602 2 8525 8568 8471 4 NOR2X1 $T=2548920 2277520 1 180 $X=2546940 $Y=2277118
X603 2 8613 8609 8608 4 NOR2X1 $T=2559480 2267440 1 180 $X=2557500 $Y=2267038
X604 2 8568 8609 8646 4 NOR2X1 $T=2572680 2267440 1 180 $X=2570700 $Y=2267038
X605 2 8685 8609 8680 4 NOR2X1 $T=2581920 2267440 1 180 $X=2579940 $Y=2267038
X606 2 8574 8313 8685 4 NOR2X1 $T=2585880 2317840 0 180 $X=2583900 $Y=2312400
X607 48 47 4 2 1785 NOR2X2 $T=770220 2247280 1 0 $X=770218 $Y=2241840
X608 81 2411 4 2 2503 NOR2X2 $T=976140 2237200 1 0 $X=976138 $Y=2231760
X609 2049 2615 4 2 2598 NOR2X2 $T=1007160 2348080 1 180 $X=1003860 $Y=2347678
X610 1874 2671 4 2 2633 NOR2X2 $T=1011780 2368240 1 180 $X=1008480 $Y=2367838
X611 2633 2598 4 2 2653 NOR2X2 $T=1016400 2388400 1 0 $X=1016398 $Y=2382960
X612 2080 2733 4 2 2731 NOR2X2 $T=1038180 2368240 1 180 $X=1034880 $Y=2367838
X613 2808 2731 4 2 2771 NOR2X2 $T=1051380 2388400 0 180 $X=1048080 $Y=2382960
X614 1912 2957 4 2 2999 NOR2X2 $T=1101540 2378320 1 0 $X=1101538 $Y=2372880
X615 1903 3295 4 2 3326 NOR2X2 $T=1176120 2378320 1 0 $X=1176118 $Y=2372880
X616 2596 3308 4 2 3337 NOR2X2 $T=1186680 2348080 0 0 $X=1186678 $Y=2347678
X617 3326 3337 4 2 3333 NOR2X2 $T=1189980 2388400 1 180 $X=1186680 $Y=2387998
X618 2226 3497 4 2 3483 NOR2X2 $T=1219020 2348080 1 180 $X=1215720 $Y=2347678
X619 2191 3445 4 2 3517 NOR2X2 $T=1217700 2368240 0 0 $X=1217698 $Y=2367838
X620 3517 3483 4 2 3516 NOR2X2 $T=1223640 2368240 0 0 $X=1223638 $Y=2367838
X621 2445 3597 4 2 3683 NOR2X2 $T=1241460 2348080 0 0 $X=1241458 $Y=2347678
X622 2649 3694 4 2 3667 NOR2X2 $T=1255320 2327920 0 180 $X=1252020 $Y=2322480
X623 2366 3744 4 2 3766 NOR2X2 $T=1269840 2348080 0 0 $X=1269838 $Y=2347678
X624 3766 3712 4 2 3695 NOR2X2 $T=1279080 2388400 0 180 $X=1275780 $Y=2382960
X625 3917 3914 4 2 3971 NOR2X2 $T=1314720 2327920 1 0 $X=1314718 $Y=2322480
X626 4163 4165 4 2 4028 NOR2X2 $T=1374120 2388400 0 180 $X=1370820 $Y=2382960
X627 4230 4295 4 2 4273 NOR2X2 $T=1406460 2247280 0 0 $X=1406458 $Y=2246878
X628 4294 4292 4 2 4230 NOR2X2 $T=1407120 2267440 1 0 $X=1407118 $Y=2262000
X629 4733 4719 4 2 4720 NOR2X2 $T=1531860 2388400 1 0 $X=1531858 $Y=2382960
X630 4851 4854 4 2 4737 NOR2X2 $T=1545720 2327920 0 180 $X=1542420 $Y=2322480
X631 4769 4767 4 2 4719 NOR2X2 $T=1545060 2388400 0 0 $X=1545058 $Y=2387998
X632 5217 5857 4 2 5860 NOR2X2 $T=1820940 2287600 0 180 $X=1817640 $Y=2282160
X633 3331 377 4 2 6284 NOR2X2 $T=1934460 2338000 1 0 $X=1934458 $Y=2332560
X634 6314 6290 4 2 6319 NOR2X2 $T=1941060 2307760 0 180 $X=1937760 $Y=2302320
X635 3944 6410 4 2 6431 NOR2X2 $T=1959540 2257360 0 0 $X=1959538 $Y=2256958
X636 3670 394 4 2 6501 NOR2X2 $T=1981980 2368240 1 0 $X=1981978 $Y=2362800
X637 6505 6501 4 2 6473 NOR2X2 $T=1983960 2317840 1 0 $X=1983958 $Y=2312400
X638 3669 398 4 2 6505 NOR2X2 $T=1992540 2348080 0 0 $X=1992538 $Y=2347678
X639 6959 423 4 2 424 NOR2X2 $T=2107380 2237200 0 180 $X=2104080 $Y=2231760
X640 438 436 4 2 7039 NOR2X2 $T=2145000 2267440 0 180 $X=2141700 $Y=2262000
X641 7450 7352 4 2 7448 NOR2X2 $T=2253240 2267440 1 180 $X=2249940 $Y=2267038
X642 7512 7464 4 2 7482 NOR2X2 $T=2270400 2287600 0 0 $X=2270398 $Y=2287198
X643 7818 7654 4 2 7828 NOR2X2 $T=2354220 2317840 1 0 $X=2354218 $Y=2312400
X644 7828 7862 4 2 7860 NOR2X2 $T=2370720 2287600 1 180 $X=2367420 $Y=2287198
X645 7846 7847 4 2 7862 NOR2X2 $T=2369400 2317840 0 0 $X=2369398 $Y=2317438
X646 8088 8039 4 2 8122 NOR2X2 $T=2440680 2257360 0 0 $X=2440678 $Y=2256958
X647 8172 8123 4 2 8187 NOR2X2 $T=2455200 2277520 1 0 $X=2455198 $Y=2272080
X648 8186 8215 4 2 8201 NOR2X2 $T=2465100 2297680 1 180 $X=2461800 $Y=2297278
X649 65 2224 4 2 2228 OR2XL $T=901560 2257360 1 0 $X=901558 $Y=2251920
X650 1815 2904 4 2 3006 OR2XL $T=1079760 2348080 0 0 $X=1079758 $Y=2347678
X651 204 4729 4 2 258 OR2XL $T=1526580 2237200 0 0 $X=1526578 $Y=2236798
X652 5631 323 4 2 5655 OR2XL $T=1764840 2327920 0 0 $X=1764838 $Y=2327518
X653 5266 403 4 2 6602 OR2XL $T=2006400 2287600 0 0 $X=2006398 $Y=2287198
X654 6772 8418 4 2 8476 OR2XL $T=2535060 2388400 0 180 $X=2532420 $Y=2382960
X655 66 2332 2294 4 2 NAND2X2 $T=931260 2267440 1 180 $X=927960 $Y=2267038
X656 2351 73 2411 4 2 NAND2X2 $T=954360 2237200 1 180 $X=951060 $Y=2236798
X657 2049 2615 2613 4 2 NAND2X2 $T=1007820 2358160 1 180 $X=1004520 $Y=2357758
X658 1912 2957 2959 4 2 NAND2X2 $T=1096920 2378320 0 180 $X=1093620 $Y=2372880
X659 3001 1609 2998 4 2 NAND2X2 $T=1101540 2348080 0 0 $X=1101538 $Y=2347678
X660 2974 3082 3099 4 2 NAND2X2 $T=1129260 2297680 0 180 $X=1125960 $Y=2292240
X661 1903 3295 3283 4 2 NAND2X2 $T=1178100 2368240 1 180 $X=1174800 $Y=2367838
X662 3333 3516 157 4 2 NAND2X2 $T=1242120 2398480 0 180 $X=1238820 $Y=2393040
X663 4067 4087 4121 4 2 NAND2X2 $T=1364220 2327920 1 0 $X=1364218 $Y=2322480
X664 3239 216 4363 4 2 NAND2X2 $T=1431540 2388400 1 180 $X=1428240 $Y=2387998
X665 2735 220 4412 4 2 NAND2X2 $T=1441440 2388400 0 0 $X=1441438 $Y=2387998
X666 4409 232 4476 4 2 NAND2X2 $T=1460580 2388400 1 180 $X=1457280 $Y=2387998
X667 4657 4659 4294 4 2 NAND2X2 $T=1512060 2297680 1 180 $X=1508760 $Y=2297278
X668 3150 358 6002 4 2 NAND2X2 $T=1852620 2317840 0 180 $X=1849320 $Y=2312400
X669 5990 6044 6020 4 2 NAND2X2 $T=1867140 2297680 1 180 $X=1863840 $Y=2297278
X670 3896 6299 380 4 2 NAND2X2 $T=1935120 2237200 0 180 $X=1931820 $Y=2231760
X671 3379 382 6322 4 2 NAND2X2 $T=1940400 2338000 1 180 $X=1937100 $Y=2337598
X672 6473 6444 6466 4 2 NAND2X2 $T=1974720 2317840 1 0 $X=1974718 $Y=2312400
X673 3670 394 397 4 2 NAND2X2 $T=1981980 2378320 1 0 $X=1981978 $Y=2372880
X674 7450 7352 7449 4 2 NAND2X2 $T=2251260 2277520 1 180 $X=2247960 $Y=2277118
X675 7639 7574 7623 4 2 NAND2X2 $T=2302740 2297680 0 180 $X=2299440 $Y=2292240
X676 8172 8123 8199 4 2 NAND2X2 $T=2459160 2277520 1 180 $X=2455860 $Y=2277118
X677 8217 8122 8241 4 2 NAND2X2 $T=2475660 2257360 0 0 $X=2475658 $Y=2256958
X678 1785 2 1796 46 4 1643 AOI21X4 $T=778140 2267440 1 180 $X=771540 $Y=2267038
X679 1876 2 56 1799 4 1899 AOI21X4 $T=803880 2317840 1 0 $X=803878 $Y=2312400
X680 67 2 2318 2313 4 2308 AOI21X4 $T=933900 2287600 1 180 $X=927300 $Y=2287198
X681 69 2 2351 2306 4 2444 AOI21X4 $T=939180 2247280 0 0 $X=939178 $Y=2246878
X682 83 2 2454 2488 4 2522 AOI21X4 $T=975480 2267440 0 0 $X=975478 $Y=2267038
X683 2503 2 86 2521 4 2612 AOI21X4 $T=984060 2237200 1 0 $X=984058 $Y=2231760
X684 2616 2 2599 2634 4 2664 AOI21X4 $T=1006500 2398480 0 0 $X=1006498 $Y=2398078
X685 2667 2 2699 2696 4 2714 AOI21X4 $T=1027620 2277520 0 0 $X=1027618 $Y=2277118
X686 2616 2 2653 2740 4 2738 AOI21X4 $T=1045440 2398480 1 180 $X=1038840 $Y=2398078
X687 2771 2 2740 2810 4 97 AOI21X4 $T=1050720 2398480 0 0 $X=1050718 $Y=2398078
X688 3035 2 111 107 4 2978 AOI21X4 $T=1112760 2408560 0 180 $X=1106160 $Y=2403120
X689 2616 2 3047 3021 4 3106 AOI21X4 $T=1116720 2388400 1 0 $X=1116718 $Y=2382960
X690 2960 2 3082 3098 4 3092 AOI21X4 $T=1124640 2287600 1 0 $X=1124638 $Y=2282160
X691 2616 2 3101 3127 4 3121 AOI21X4 $T=1142460 2398480 1 180 $X=1135860 $Y=2398078
X692 3019 2 3292 3296 4 3299 AOI21X4 $T=1174140 2297680 1 0 $X=1174138 $Y=2292240
X693 3971 2 180 3980 4 4069 AOI21X4 $T=1331220 2317840 0 0 $X=1331218 $Y=2317438
X694 4273 2 200 4233 4 4101 AOI21X4 $T=1402500 2247280 1 180 $X=1395900 $Y=2246878
X695 4122 2 4379 4362 4 4396 AOI21X4 $T=1434180 2368240 1 0 $X=1434178 $Y=2362800
X696 4420 2 4409 4461 4 4472 AOI21X4 $T=1448700 2368240 0 0 $X=1448698 $Y=2367838
X697 4461 2 232 4491 4 4502 AOI21X4 $T=1459920 2378320 1 0 $X=1459918 $Y=2372880
X698 248 2 4720 255 4 254 AOI21X4 $T=1527900 2408560 1 180 $X=1521300 $Y=2408158
X699 4501 2 5860 5907 4 5916 AOI21X4 $T=1825560 2287600 1 0 $X=1825558 $Y=2282160
X700 6023 2 5990 6040 4 6077 AOI21X4 $T=1863180 2277520 1 0 $X=1863178 $Y=2272080
X701 6044 2 6040 6078 4 6037 AOI21X4 $T=1873740 2297680 1 0 $X=1873738 $Y=2292240
X702 6041 2 6319 6348 4 6461 AOI21X4 $T=1941060 2297680 0 0 $X=1941058 $Y=2297278
X703 6803 2 6761 6817 4 6821 AOI21X4 $T=2068440 2267440 1 0 $X=2068438 $Y=2262000
X704 6946 2 6948 6961 4 6962 AOI21X4 $T=2102760 2368240 1 0 $X=2102758 $Y=2362800
X705 7484 2 7319 7498 4 7636 AOI21X4 $T=2262480 2267440 1 0 $X=2262478 $Y=2262000
X706 7626 2 7643 7671 4 7673 AOI21X4 $T=2312640 2257360 0 0 $X=2312638 $Y=2256958
X707 7786 2 7860 7863 4 7879 AOI21X4 $T=2366760 2277520 0 0 $X=2366758 $Y=2277118
X708 8089 2 8217 8249 4 8254 AOI21X4 $T=2471700 2267440 0 0 $X=2471698 $Y=2267038
X709 1783 2 1785 4 1641 AND2X2 $T=773520 2297680 1 180 $X=770880 $Y=2297278
X710 1783 2 1827 4 1900 AND2X2 $T=788040 2267440 1 0 $X=788038 $Y=2262000
X711 2189 2 2176 4 2196 AND2X2 $T=896280 2327920 0 0 $X=896278 $Y=2327518
X712 2318 2 2294 4 2368 AND2X2 $T=939840 2287600 0 0 $X=939838 $Y=2287198
X713 2454 2 78 4 2482 AND2X2 $T=965580 2277520 1 0 $X=965578 $Y=2272080
X714 2599 2 2613 4 2614 AND2X2 $T=1003860 2388400 1 0 $X=1003858 $Y=2382960
X715 3283 2 3317 4 3271 AND2X2 $T=1173480 2398480 1 180 $X=1170840 $Y=2398078
X716 3632 2 3594 4 3595 AND2X2 $T=1242780 2287600 1 180 $X=1240140 $Y=2287198
X717 3883 2 3898 4 3913 AND2X2 $T=1306800 2267440 1 0 $X=1306798 $Y=2262000
X718 3993 2 3972 4 3958 AND2X2 $T=1335840 2338000 1 180 $X=1333200 $Y=2337598
X719 4066 2 4086 4 4087 AND2X2 $T=1356960 2307760 0 0 $X=1356958 $Y=2307358
X720 4085 2 4086 4 4117 AND2X2 $T=1357620 2287600 1 0 $X=1357618 $Y=2282160
X721 4409 2 4412 4 4399 AND2X2 $T=1442760 2378320 1 180 $X=1440120 $Y=2377918
X722 4720 2 257 4 261 AND2X2 $T=1533180 2408560 0 0 $X=1533178 $Y=2408158
X723 277 2 281 4 4952 AND2X2 $T=1591920 2237200 0 180 $X=1589280 $Y=2231760
X724 5102 2 5105 4 5106 AND2X2 $T=1623600 2277520 0 0 $X=1623598 $Y=2277118
X725 5151 2 5219 4 302 AND2X2 $T=1657920 2398480 0 0 $X=1657918 $Y=2398078
X726 328 2 319 4 5488 AND2X2 $T=1731180 2287600 0 180 $X=1728540 $Y=2282160
X727 5594 2 329 4 5627 AND2X2 $T=1754280 2358160 1 0 $X=1754278 $Y=2352720
X728 5655 2 5713 4 5708 AND2X2 $T=1793220 2338000 0 180 $X=1790580 $Y=2332560
X729 5655 2 5724 4 5757 AND2X2 $T=1793220 2338000 0 0 $X=1793218 $Y=2337598
X730 5891 2 350 4 5877 AND2X2 $T=1826880 2388400 0 180 $X=1824240 $Y=2382960
X731 5990 2 6002 4 6006 AND2X2 $T=1856580 2277520 1 0 $X=1856578 $Y=2272080
X732 6222 2 6075 4 6235 AND2X2 $T=1915320 2398480 0 0 $X=1915318 $Y=2398078
X733 3331 2 377 4 6234 AND2X2 $T=1924560 2338000 0 180 $X=1921920 $Y=2332560
X734 375 2 6134 4 6253 AND2X2 $T=1929180 2378320 0 180 $X=1926540 $Y=2372880
X735 6789 2 6730 4 6817 AND2X2 $T=2070420 2257360 0 0 $X=2070418 $Y=2256958
X736 6855 2 6853 4 418 AND2X2 $T=2083620 2408560 1 180 $X=2080980 $Y=2408158
X737 7643 2 7623 4 7625 AND2X2 $T=2307360 2257360 1 180 $X=2304720 $Y=2256958
X738 8099 2 8009 4 475 AND2X2 $T=2430120 2237200 1 180 $X=2427480 $Y=2236798
X739 1611 4 1623 2 1556 NAND2X4 $T=724020 2338000 0 0 $X=724018 $Y=2337598
X740 2691 4 2651 2 2740 NAND2X4 $T=1035540 2398480 1 0 $X=1035538 $Y=2393040
X741 2771 4 2653 2 99 NAND2X4 $T=1061280 2398480 0 0 $X=1061278 $Y=2398078
X742 4124 4 4121 2 4122 NAND2X4 $T=1369500 2327920 1 180 $X=1364880 $Y=2327518
X743 288 4 2880 2 5168 NAND2X4 $T=1610400 2287600 1 0 $X=1610398 $Y=2282160
X744 369 4 3159 2 6191 NAND2X4 $T=1898160 2317840 0 0 $X=1898158 $Y=2317438
X745 6189 4 6260 2 6290 NAND2X4 $T=1931820 2307760 0 180 $X=1927200 $Y=2302320
X746 1687 1642 4 2 1623 OR2X2 $T=736560 2338000 1 180 $X=733920 $Y=2337598
X747 2104 2168 4 2 2176 OR2X2 $T=892320 2307760 1 0 $X=892318 $Y=2302320
X748 2350 2352 4 2 2353 OR2X2 $T=939840 2327920 1 0 $X=939838 $Y=2322480
X749 2436 43 4 2 2356 OR2X2 $T=961620 2327920 0 180 $X=958980 $Y=2322480
X750 2260 82 4 2 2500 OR2X2 $T=976140 2307760 0 0 $X=976138 $Y=2307358
X751 2262 82 4 2 2520 OR2X2 $T=982740 2307760 0 0 $X=982738 $Y=2307358
X752 2714 2689 4 2 2718 OR2X2 $T=1030920 2317840 1 0 $X=1030918 $Y=2312400
X753 2751 2731 4 2 2770 OR2X2 $T=1042800 2388400 1 0 $X=1042798 $Y=2382960
X754 3099 3146 4 2 3205 OR2X2 $T=1147740 2287600 0 0 $X=1147738 $Y=2287198
X755 3742 3800 4 2 3807 OR2X2 $T=1287000 2257360 1 0 $X=1286998 $Y=2251920
X756 4278 206 4 2 4274 OR2X2 $T=1413060 2358160 0 180 $X=1410420 $Y=2352720
X757 4328 4318 4 2 4305 OR2X2 $T=1416360 2338000 1 180 $X=1413720 $Y=2337598
X758 4678 4676 4 2 4659 OR2X2 $T=1514700 2317840 0 180 $X=1512060 $Y=2312400
X759 4711 4707 4 2 4678 OR2X2 $T=1523940 2307760 1 180 $X=1521300 $Y=2307358
X760 4886 4902 4 2 4776 OR2X2 $T=1570140 2257360 1 180 $X=1567500 $Y=2256958
X761 5032 279 4 2 5030 OR2X2 $T=1602480 2257360 0 180 $X=1599840 $Y=2251920
X762 5082 5046 4 2 5118 OR2X2 $T=1618320 2368240 1 0 $X=1618318 $Y=2362800
X763 279 281 4 2 5157 OR2X2 $T=1631520 2247280 1 0 $X=1631518 $Y=2241840
X764 5170 5159 4 2 5151 OR2X2 $T=1642080 2388400 1 180 $X=1639440 $Y=2387998
X765 298 299 4 2 5219 OR2X2 $T=1644720 2398480 0 0 $X=1644718 $Y=2398078
X766 273 5157 4 2 5230 OR2X2 $T=1645380 2257360 1 0 $X=1645378 $Y=2251920
X767 277 5230 4 2 5231 OR2X2 $T=1657260 2267440 1 0 $X=1657258 $Y=2262000
X768 5328 309 4 2 5341 OR2X2 $T=1691580 2408560 1 0 $X=1691578 $Y=2403120
X769 271 5482 4 2 5628 OR2X2 $T=1756920 2378320 1 0 $X=1756918 $Y=2372880
X770 275 5628 4 2 5648 OR2X2 $T=1764840 2398480 1 0 $X=1764838 $Y=2393040
X771 260 5648 4 2 5651 OR2X2 $T=1772760 2398480 0 180 $X=1770120 $Y=2393040
X772 348 5924 4 2 6014 OR2X2 $T=1840740 2388400 1 0 $X=1840738 $Y=2382960
X773 321 6014 4 2 6062 OR2X2 $T=1861200 2388400 1 0 $X=1861198 $Y=2382960
X774 362 6062 4 2 363 OR2X2 $T=1874400 2408560 1 0 $X=1874398 $Y=2403120
X775 3896 6299 4 2 379 OR2X2 $T=1930500 2247280 1 0 $X=1930498 $Y=2241840
X776 6431 6442 4 2 6440 OR2X2 $T=1970100 2257360 0 180 $X=1967460 $Y=2251920
X777 338 5897 4 2 6647 OR2X2 $T=2013660 2388400 0 0 $X=2013658 $Y=2387998
X778 6662 6648 4 2 6652 OR2X2 $T=2028840 2297680 0 180 $X=2026200 $Y=2292240
X779 342 6647 4 2 6678 OR2X2 $T=2028180 2398480 0 0 $X=2028178 $Y=2398078
X780 6789 6730 4 2 6803 OR2X2 $T=2070420 2247280 0 0 $X=2070418 $Y=2246878
X781 6855 6853 4 2 425 OR2X2 $T=2086260 2408560 0 0 $X=2086258 $Y=2408158
X782 6866 6867 4 2 6948 OR2X2 $T=2087580 2368240 1 0 $X=2087578 $Y=2362800
X783 6870 6804 4 2 6864 OR2X2 $T=2090220 2327920 1 180 $X=2087580 $Y=2327518
X784 7011 7006 4 2 435 OR2X2 $T=2128500 2408560 1 180 $X=2125860 $Y=2408158
X785 7167 7185 4 2 7202 OR2X2 $T=2181960 2287600 1 0 $X=2181958 $Y=2282160
X786 8467 8450 4 2 8475 OR2X2 $T=2528460 2307760 0 180 $X=2525820 $Y=2302320
X787 8461 501 4 2 8473 OR2X2 $T=2533740 2277520 0 180 $X=2531100 $Y=2272080
X788 8549 8546 4 2 8569 OR2X2 $T=2544300 2327920 1 0 $X=2544298 $Y=2322480
X789 8613 8612 4 2 8634 OR2X2 $T=2564760 2277520 0 0 $X=2564758 $Y=2277118
X790 8611 8556 4 2 8648 OR2X2 $T=2567400 2338000 0 0 $X=2567398 $Y=2337598
X791 1827 4 2 54 1873 NAND2XL $T=797280 2257360 1 0 $X=797278 $Y=2251920
X792 2145 4 2 2176 2136 NAND2XL $T=888360 2327920 1 180 $X=886380 $Y=2327518
X793 2196 4 2 2174 2262 NAND2XL $T=899580 2327920 1 0 $X=899578 $Y=2322480
X794 2380 4 2 2353 2439 NAND2XL $T=949080 2348080 1 0 $X=949078 $Y=2342640
X795 2438 4 2 2356 2426 NAND2XL $T=962940 2338000 0 180 $X=960960 $Y=2332560
X796 43 4 2 2436 2438 NAND2XL $T=969540 2327920 0 180 $X=967560 $Y=2322480
X797 3152 4 2 3139 3102 NAND2XL $T=1141800 2307760 0 180 $X=1139820 $Y=2302320
X798 128 4 2 127 3204 NAND2XL $T=1168200 2237200 0 180 $X=1166220 $Y=2231760
X799 147 4 2 148 3494 NAND2XL $T=1213080 2237200 1 0 $X=1213078 $Y=2231760
X800 3666 4 2 3672 3685 NAND2XL $T=1254000 2277520 0 0 $X=1253998 $Y=2277118
X801 3694 4 2 2649 3706 NAND2XL $T=1259940 2327920 1 0 $X=1259938 $Y=2322480
X802 3751 4 2 3526 3753 NAND2XL $T=1275780 2257360 0 0 $X=1275778 $Y=2256958
X803 3764 4 2 3788 3809 NAND2XL $T=1283700 2398480 1 0 $X=1283698 $Y=2393040
X804 3794 4 2 2648 3881 NAND2XL $T=1292940 2287600 0 0 $X=1292938 $Y=2287198
X805 195 4 2 192 4143 NAND2XL $T=1386000 2317840 0 0 $X=1385998 $Y=2317438
X806 201 4 2 196 4219 NAND2XL $T=1387980 2277520 0 180 $X=1386000 $Y=2272080
X807 209 4 2 4314 4220 NAND2XL $T=1413720 2327920 0 180 $X=1411740 $Y=2322480
X808 4330 4 2 4305 4291 NAND2XL $T=1413720 2368240 0 180 $X=1411740 $Y=2362800
X809 5151 4 2 5069 5137 NAND2XL $T=1635480 2398480 1 180 $X=1633500 $Y=2398078
X810 5220 4 2 5151 5249 NAND2XL $T=1655280 2388400 0 0 $X=1655278 $Y=2387998
X811 5159 4 2 5170 5220 NAND2XL $T=1657920 2388400 1 0 $X=1657918 $Y=2382960
X812 309 4 2 5283 5258 NAND2XL $T=1678380 2408560 0 180 $X=1676400 $Y=2403120
X813 5313 4 2 5312 310 NAND2XL $T=1686960 2358160 0 180 $X=1684980 $Y=2352720
X814 323 4 2 5631 5724 NAND2XL $T=1772760 2327920 0 0 $X=1772758 $Y=2327518
X815 339 4 2 316 5707 NAND2XL $T=1782000 2297680 0 0 $X=1781998 $Y=2297278
X816 5150 4 2 329 5754 NAND2XL $T=1805760 2317840 1 0 $X=1805758 $Y=2312400
X817 365 4 2 5645 6133 NAND2XL $T=1882980 2368240 1 0 $X=1882978 $Y=2362800
X818 6142 4 2 375 6239 NAND2XL $T=1919940 2388400 0 0 $X=1919938 $Y=2387998
X819 375 4 2 6269 6305 NAND2XL $T=1939740 2368240 1 180 $X=1937760 $Y=2367838
X820 6267 4 2 375 6397 NAND2XL $T=1947000 2368240 0 0 $X=1946998 $Y=2367838
X821 403 4 2 5266 6619 NAND2XL $T=2018280 2277520 1 180 $X=2016300 $Y=2277118
X822 6137 4 2 6709 6805 NAND2XL $T=2063160 2327920 1 0 $X=2063158 $Y=2322480
X823 6858 4 2 6864 6892 NAND2XL $T=2093520 2307760 1 0 $X=2093518 $Y=2302320
X824 7075 4 2 6042 7182 NAND2XL $T=2171400 2408560 1 0 $X=2171398 $Y=2403120
X825 7075 4 2 7179 7181 NAND2XL $T=2181300 2398480 1 180 $X=2179320 $Y=2398078
X826 6042 4 2 7179 7184 NAND2XL $T=2189220 2408560 1 180 $X=2187240 $Y=2408158
X827 8086 4 2 8082 8173 NAND2XL $T=2450580 2338000 0 0 $X=2450578 $Y=2337598
X828 8199 4 2 8176 484 NAND2XL $T=2460480 2237200 0 0 $X=2460478 $Y=2236798
X829 7719 4 2 472 8472 NAND2XL $T=2528460 2297680 1 0 $X=2528458 $Y=2292240
X830 7719 4 2 8424 505 NAND2XL $T=2533740 2287600 0 0 $X=2533738 $Y=2287198
X831 8418 4 2 6772 8505 NAND2XL $T=2537700 2378320 1 0 $X=2537698 $Y=2372880
X832 8577 4 2 8569 8632 NAND2XL $T=2560140 2307760 0 0 $X=2560138 $Y=2307358
X833 8615 4 2 8648 8668 NAND2XL $T=2572020 2307760 0 0 $X=2572018 $Y=2307358
X834 8729 4 2 8666 8714 NAND2XL $T=2593800 2287600 1 180 $X=2591820 $Y=2287198
X835 2756 3023 4 2 INVX4 $T=1084380 2307760 0 0 $X=1084378 $Y=2307358
X836 97 3035 4 2 INVX4 $T=1118700 2408560 1 0 $X=1118698 $Y=2403120
X837 4069 4067 4 2 INVX4 $T=1354320 2327920 0 180 $X=1351680 $Y=2322480
X838 238 231 4 2 INVX4 $T=1485660 2247280 1 180 $X=1483020 $Y=2246878
X839 4746 248 4 2 INVX4 $T=1537140 2348080 1 180 $X=1534500 $Y=2347678
X840 291 281 4 2 INVX4 $T=1619640 2237200 1 0 $X=1619638 $Y=2231760
X841 4501 5909 4 2 INVX4 $T=1830180 2277520 0 0 $X=1830178 $Y=2277118
X842 5714 6042 4 2 INVX4 $T=1861200 2398480 1 0 $X=1861198 $Y=2393040
X843 5633 6737 4 2 INVX4 $T=2049960 2368240 1 0 $X=2049958 $Y=2362800
X844 5280 6736 4 2 INVX4 $T=2061840 2358160 0 0 $X=2061838 $Y=2357758
X845 7636 7626 4 2 INVX4 $T=2306040 2267440 1 180 $X=2303400 $Y=2267038
X846 7786 7794 4 2 INVX4 $T=2350920 2277520 0 180 $X=2348280 $Y=2272080
X847 7879 478 4 2 INVX4 $T=2442000 2257360 1 0 $X=2441998 $Y=2251920
X848 1737 1593 2 1733 1734 4 AOI21X1 $T=759000 2317840 0 180 $X=756360 $Y=2312400
X849 1638 1756 2 1593 1752 4 AOI21X1 $T=762960 2327920 0 180 $X=760320 $Y=2322480
X850 1724 1756 2 1723 1755 4 AOI21X1 $T=762960 2338000 0 180 $X=760320 $Y=2332560
X851 1796 1827 2 1849 1898 4 AOI21X1 $T=797280 2257360 0 0 $X=797278 $Y=2256958
X852 2176 2106 2 2151 2225 4 AOI21X1 $T=900240 2338000 1 0 $X=900238 $Y=2332560
X853 2353 2343 2 2346 2344 4 AOI21X1 $T=941160 2358160 0 180 $X=938520 $Y=2352720
X854 2346 2356 2 2354 2310 4 AOI21X1 $T=943140 2338000 0 180 $X=940500 $Y=2332560
X855 2974 2756 2 2960 2958 4 AOI21X1 $T=1098240 2287600 1 180 $X=1095600 $Y=2287198
X856 3139 3198 2 3160 3158 4 AOI21X1 $T=1150380 2307760 0 180 $X=1147740 $Y=2302320
X857 3218 3198 2 3243 3244 4 AOI21X1 $T=1162920 2297680 0 0 $X=1162918 $Y=2297278
X858 3243 3220 2 3255 3294 4 AOI21X1 $T=1165560 2277520 0 0 $X=1165558 $Y=2277118
X859 3258 3198 2 3274 3275 4 AOI21X1 $T=1170840 2297680 0 0 $X=1170838 $Y=2297278
X860 3425 3328 2 3430 3431 4 AOI21X1 $T=1203840 2388400 1 0 $X=1203838 $Y=2382960
X861 3592 132 2 3518 3566 4 AOI21X1 $T=1234860 2408560 0 180 $X=1232220 $Y=2403120
X862 166 3728 2 3749 3745 4 AOI21X1 $T=1275780 2398480 1 180 $X=1273140 $Y=2398078
X863 3695 166 2 3720 3827 4 AOI21X1 $T=1290960 2398480 0 0 $X=1290958 $Y=2398078
X864 3788 166 2 3811 173 4 AOI21X1 $T=1296240 2398480 0 0 $X=1296238 $Y=2398078
X865 132 3886 2 3853 3899 4 AOI21X1 $T=1306800 2408560 1 0 $X=1306798 $Y=2403120
X866 3913 177 2 3946 3970 4 AOI21X1 $T=1329240 2267440 1 0 $X=1329238 $Y=2262000
X867 4212 4214 2 4216 4221 4 AOI21X1 $T=1393920 2338000 0 0 $X=1393918 $Y=2337598
X868 4274 4272 2 4276 4281 4 AOI21X1 $T=1401180 2378320 1 0 $X=1401178 $Y=2372880
X869 4305 4276 2 4343 4309 4 AOI21X1 $T=1419660 2378320 1 0 $X=1419658 $Y=2372880
X870 4660 248 2 4655 4643 4 AOI21X1 $T=1511400 2388400 0 180 $X=1508760 $Y=2382960
X871 284 5030 2 5031 267 4 AOI21X1 $T=1603140 2237200 1 0 $X=1603138 $Y=2231760
X872 302 293 2 5258 5265 4 AOI21X1 $T=1665180 2408560 1 0 $X=1665178 $Y=2403120
X873 5069 5264 2 293 5260 4 AOI21X1 $T=1670460 2388400 0 180 $X=1667820 $Y=2382960
X874 5426 5439 2 5441 5340 4 AOI21X1 $T=1714680 2388400 0 0 $X=1714678 $Y=2387998
X875 5501 5593 2 5606 5673 4 AOI21X1 $T=1755600 2257360 1 0 $X=1755598 $Y=2251920
X876 6120 6116 2 6102 6112 4 AOI21X1 $T=1890240 2358160 1 180 $X=1887600 $Y=2357758
X877 6142 370 2 6120 6192 4 AOI21X1 $T=1906080 2388400 1 180 $X=1903440 $Y=2387998
X878 6621 6652 2 6650 6692 4 AOI21X1 $T=2024880 2287600 0 0 $X=2024878 $Y=2287198
X879 425 427 2 418 7012 4 AOI21X1 $T=2112660 2408560 0 0 $X=2112658 $Y=2408158
X880 7202 7200 2 7229 7282 4 AOI21X1 $T=2193840 2257360 0 0 $X=2193838 $Y=2256958
X881 7229 7284 2 7304 7317 4 AOI21X1 $T=2212320 2267440 1 0 $X=2212318 $Y=2262000
X882 8357 8471 2 8519 503 4 AOI21X1 $T=2545620 2267440 1 180 $X=2542980 $Y=2267038
X883 8463 493 2 8357 8596 4 AOI21X1 $T=2544300 2267440 1 0 $X=2544298 $Y=2262000
X884 8608 493 2 8599 8598 4 AOI21X1 $T=2557500 2267440 0 180 $X=2554860 $Y=2262000
X885 8569 8618 2 8516 8614 4 AOI21X1 $T=2561460 2297680 1 180 $X=2558820 $Y=2297278
X886 8646 493 2 8645 8643 4 AOI21X1 $T=2571360 2267440 0 180 $X=2568720 $Y=2262000
X887 8648 8649 2 8647 8528 4 AOI21X1 $T=2572680 2297680 1 180 $X=2570040 $Y=2297278
X888 8680 493 2 8681 8679 4 AOI21X1 $T=2578620 2267440 1 0 $X=2578618 $Y=2262000
X889 1787 1687 4 1752 2 1786 OAI21X2 $T=773520 2338000 1 0 $X=773518 $Y=2332560
X890 51 1687 4 52 2 1848 OAI21X2 $T=798600 2338000 1 180 $X=793320 $Y=2337598
X891 1871 1687 4 1847 2 1886 OAI21X2 $T=801240 2297680 1 180 $X=795960 $Y=2297278
X892 2105 1899 4 2088 2 2102 OAI21X2 $T=869220 2348080 0 180 $X=863940 $Y=2342640
X893 2148 1899 4 2167 2 2146 OAI21X2 $T=887040 2348080 0 0 $X=887038 $Y=2347678
X894 2294 2242 4 2259 2 2306 OAI21X2 $T=927960 2257360 0 180 $X=922680 $Y=2251920
X895 2411 80 4 2444 2 2521 OAI21X2 $T=969540 2237200 1 180 $X=964260 $Y=2236798
X896 2747 2808 4 2769 2 2810 OAI21X2 $T=1053360 2358160 1 180 $X=1048080 $Y=2357758
X897 2842 2919 4 2920 2 2960 OAI21X2 $T=1082400 2287600 1 0 $X=1082398 $Y=2282160
X898 2998 2905 4 3004 2 109 OAI21X2 $T=1100220 2358160 0 0 $X=1100218 $Y=2357758
X899 3022 3023 4 3011 2 3026 OAI21X2 $T=1110780 2307760 0 180 $X=1105500 $Y=2302320
X900 2980 2978 4 2998 2 3039 OAI21X2 $T=1113420 2368240 0 180 $X=1108140 $Y=2362800
X901 3205 3023 4 3158 2 3199 OAI21X2 $T=1150380 2317840 0 180 $X=1145100 $Y=2312400
X902 3897 3917 4 3972 2 3980 OAI21X2 $T=1335840 2327920 1 180 $X=1330560 $Y=2327518
X903 4208 4230 4 4210 2 4233 OAI21X2 $T=1398540 2257360 0 0 $X=1398538 $Y=2256958
X904 250 4654 4 4642 2 200 OAI21X2 $T=1512720 2247280 0 180 $X=1507440 $Y=2241840
X905 4656 4719 4 4688 2 255 OAI21X2 $T=1527240 2388400 1 180 $X=1521960 $Y=2387998
X906 4779 4764 4 4793 2 4755 OAI21X2 $T=1539780 2287600 1 0 $X=1539778 $Y=2282160
X907 5217 5909 4 5168 2 5989 OAI21X2 $T=1832820 2257360 0 0 $X=1832818 $Y=2256958
X908 5168 5857 4 5927 2 5907 OAI21X2 $T=1835460 2287600 1 0 $X=1835458 $Y=2282160
X909 397 6505 4 6534 2 6509 OAI21X2 $T=1989900 2327920 0 0 $X=1989898 $Y=2327518
X910 6442 387 4 6409 2 6633 OAI21X2 $T=2001120 2237200 1 180 $X=1995840 $Y=2236798
X911 7862 7819 4 7859 2 7863 OAI21X2 $T=2371380 2307760 0 180 $X=2366100 $Y=2302320
X912 1555 1556 1609 4 2 XNOR2X4 $T=705540 2338000 0 0 $X=705538 $Y=2337598
X913 1735 1786 1815 4 2 XNOR2X4 $T=772200 2348080 1 0 $X=772198 $Y=2342640
X914 45 1885 1912 4 2 XNOR2X4 $T=804540 2257360 1 0 $X=804538 $Y=2251920
X915 1838 1848 2080 4 2 XNOR2X4 $T=804540 2338000 0 0 $X=804538 $Y=2337598
X916 2090 2102 2191 4 2 XNOR2X4 $T=867240 2368240 0 0 $X=867238 $Y=2367838
X917 2136 2146 2226 4 2 XNOR2X4 $T=884400 2358160 1 0 $X=884398 $Y=2352720
X918 3002 3121 3150 4 2 XNOR2X4 $T=1133220 2398480 1 0 $X=1133218 $Y=2393040
X919 3202 3199 2904 4 2 XNOR2X4 $T=1153020 2327920 1 180 $X=1141800 $Y=2327518
X920 3271 131 3331 4 2 XNOR2X4 $T=1177440 2408560 1 0 $X=1177438 $Y=2403120
X921 5985 5989 359 4 2 XNOR2X4 $T=1849980 2237200 1 0 $X=1849978 $Y=2231760
X922 7861 7831 469 4 2 XNOR2X4 $T=2368080 2277520 1 0 $X=2368078 $Y=2272080
X923 52 4 50 49 2 1796 OAI21X4 $T=791340 2257360 0 180 $X=784080 $Y=2251920
X924 1850 4 1687 1840 2 1874 OAI21X4 $T=795960 2358160 1 0 $X=795958 $Y=2352720
X925 94 4 2755 2737 2 2756 OAI21X4 $T=1046760 2287600 1 180 $X=1039500 $Y=2287198
X926 2908 4 2959 2907 2 107 OAI21X4 $T=1097580 2398480 1 180 $X=1090320 $Y=2398078
X927 4476 4 4396 4502 2 4501 OAI21X4 $T=1461900 2368240 1 0 $X=1461898 $Y=2362800
X928 6020 4 5916 6037 2 6041 OAI21X4 $T=1861860 2287600 0 0 $X=1861858 $Y=2287198
X929 6151 4 6262 6191 2 6265 OAI21X4 $T=1925220 2287600 0 180 $X=1917960 $Y=2282160
X930 6262 4 6290 6289 2 6301 OAI21X4 $T=1935120 2297680 0 180 $X=1927860 $Y=2292240
X931 6314 4 6289 6322 2 6348 OAI21X4 $T=1939740 2317840 0 0 $X=1939738 $Y=2317438
X932 6466 4 6464 6472 2 390 OAI21X4 $T=1971420 2307760 1 0 $X=1971418 $Y=2302320
X933 6821 4 6885 6897 2 6946 OAI21X4 $T=2092200 2317840 1 0 $X=2092198 $Y=2312400
X934 6992 4 426 7007 2 7009 OAI21X4 $T=2117940 2267440 0 0 $X=2117938 $Y=2267038
X935 7286 4 446 7317 2 7319 OAI21X4 $T=2212320 2257360 0 0 $X=2212318 $Y=2256958
X936 7448 4 7381 7449 2 7511 OAI21X4 $T=2257860 2257360 1 0 $X=2257858 $Y=2251920
X937 7675 4 7636 7689 2 7786 OAI21X4 $T=2328480 2277520 1 0 $X=2328478 $Y=2272080
X938 7828 4 7794 7819 2 7831 OAI21X4 $T=2361480 2277520 1 180 $X=2354220 $Y=2277118
X939 7879 4 8241 8254 2 493 OAI21X4 $T=2473680 2257360 1 0 $X=2473678 $Y=2251920
X940 5677 4 5709 2 CLKBUFX8 $T=1777380 2378320 0 0 $X=1777378 $Y=2377918
X941 6074 4 6786 2 CLKBUFX8 $T=2057880 2378320 0 0 $X=2057878 $Y=2377918
X942 2190 1899 2 4 2596 XOR2X2 $T=975480 2348080 0 0 $X=975478 $Y=2347678
X943 40 2519 2 4 2649 XOR2X2 $T=988680 2317840 0 0 $X=988678 $Y=2317438
X944 2695 2687 2 4 2224 XOR2X2 $T=1028940 2247280 1 180 $X=1022340 $Y=2246878
X945 2614 2616 2 4 3239 XOR2X2 $T=1150380 2388400 0 0 $X=1150378 $Y=2387998
X946 3809 3709 2 4 3931 XOR2X2 $T=1290300 2398480 1 0 $X=1290298 $Y=2393040
X947 3916 3928 2 4 3944 XOR2X2 $T=1315380 2257360 1 0 $X=1315378 $Y=2251920
X948 4008 4009 2 4 181 XOR2X2 $T=1345740 2368240 1 180 $X=1339140 $Y=2367838
X949 4162 4160 2 4 199 XOR2X2 $T=1378080 2287600 0 0 $X=1378078 $Y=2287198
X950 4644 4643 2 4 4165 XOR2X2 $T=1504800 2388400 0 180 $X=1498200 $Y=2382960
X951 265 5444 2 4 5508 XOR2X2 $T=1725240 2317840 0 0 $X=1725238 $Y=2317438
X952 5832 5348 2 4 344 XOR2X2 $T=1807080 2378320 1 0 $X=1807078 $Y=2372880
X953 5906 5909 2 4 366 XOR2X2 $T=1829520 2237200 0 0 $X=1829518 $Y=2236798
X954 311 5507 2 4 5942 XOR2X2 $T=1836120 2368240 0 0 $X=1836118 $Y=2367838
X955 321 6014 2 4 6059 XOR2X2 $T=1859220 2368240 0 0 $X=1859218 $Y=2367838
X956 6892 6884 2 4 421 XOR2X2 $T=2096160 2287600 0 180 $X=2089560 $Y=2282160
X957 7066 7053 2 4 437 XOR2X2 $T=2140380 2237200 1 0 $X=2140378 $Y=2231760
X958 7706 7673 2 4 462 XOR2X2 $T=2326500 2257360 0 0 $X=2326498 $Y=2256958
X959 8578 8598 2 4 511 XOR2X2 $T=2552880 2247280 0 0 $X=2552878 $Y=2246878
X960 8632 8643 2 4 514 XOR2X2 $T=2565420 2247280 0 0 $X=2565418 $Y=2246878
X961 8668 8679 2 4 519 XOR2X2 $T=2576640 2257360 1 0 $X=2576638 $Y=2251920
X962 8714 8596 2 4 525 XOR2X2 $T=2589180 2247280 0 0 $X=2589178 $Y=2246878
X963 2978 4 3021 2 INVX2 $T=1098240 2388400 1 0 $X=1098238 $Y=2382960
X964 3024 4 3047 2 INVX2 $T=1108800 2388400 1 0 $X=1108798 $Y=2382960
X965 5916 4 6023 2 INVX2 $T=1861860 2267440 0 0 $X=1861858 $Y=2267038
X966 446 4 7200 2 INVX2 $T=2182620 2257360 0 180 $X=2180640 $Y=2251920
X967 6059 4 7316 2 INVX2 $T=2215620 2358160 0 0 $X=2215618 $Y=2357758
X968 6786 4 7336 2 INVX2 $T=2291520 2338000 0 0 $X=2291518 $Y=2337598
X969 472 4 7849 2 INVX2 $T=2404380 2327920 1 0 $X=2404378 $Y=2322480
X970 6772 4 7719 2 INVX2 $T=2500740 2327920 0 0 $X=2500738 $Y=2327518
X971 1572 2 4 1608 INVXL $T=718080 2327920 1 0 $X=718078 $Y=2322480
X972 48 2 4 1827 INVXL $T=779460 2247280 0 0 $X=779458 $Y=2246878
X973 54 2 4 1849 INVXL $T=796620 2247280 1 0 $X=796618 $Y=2241840
X974 2613 2 4 2634 INVXL $T=1007160 2398480 1 0 $X=1007158 $Y=2393040
X975 3003 2 4 3020 INVXL $T=1103520 2277520 0 0 $X=1103518 $Y=2277118
X976 2980 2 4 3038 INVXL $T=1112760 2348080 1 0 $X=1112758 $Y=2342640
X977 3152 2 4 3160 INVXL $T=1144440 2307760 1 0 $X=1144438 $Y=2302320
X978 3146 2 4 3139 INVXL $T=1146420 2297680 0 180 $X=1145100 $Y=2292240
X979 3243 2 4 3309 INVXL $T=1176780 2297680 0 0 $X=1176778 $Y=2297278
X980 3611 2 4 3594 INVXL $T=1243440 2267440 1 180 $X=1242120 $Y=2267038
X981 3764 2 4 3811 INVXL $T=1288320 2398480 0 0 $X=1288318 $Y=2398078
X982 4221 2 4 4272 INVXL $T=1397880 2378320 1 0 $X=1397878 $Y=2372880
X983 4656 2 4 4655 INVXL $T=1510080 2388400 1 180 $X=1508760 $Y=2387998
X984 4745 2 4 4707 INVXL $T=1533840 2307760 0 180 $X=1532520 $Y=2302320
X985 5676 2 4 5689 INVXL $T=1777380 2338000 1 0 $X=1777378 $Y=2332560
X986 5724 2 4 5716 INVXL $T=1785300 2338000 1 180 $X=1783980 $Y=2337598
X987 342 2 4 340 INVXL $T=1800480 2378320 0 0 $X=1800478 $Y=2377918
X988 336 2 4 354 INVXL $T=1836120 2338000 0 0 $X=1836118 $Y=2337598
X989 8009 2 4 8103 INVXL $T=2434740 2247280 1 0 $X=2434738 $Y=2241840
X990 158 159 3627 2 3625 3671 4 AOI31X1 $T=1246740 2237200 1 0 $X=1246738 $Y=2231760
X991 1685 1757 2 4 1903 XNOR2X2 $T=760980 2358160 0 0 $X=760978 $Y=2357758
X992 1626 1818 2 4 1902 XNOR2X2 $T=782100 2338000 1 0 $X=782098 $Y=2332560
X993 1873 1886 2 4 1913 XNOR2X2 $T=807840 2297680 0 0 $X=807838 $Y=2297278
X994 60 61 2 4 2049 XNOR2X2 $T=832920 2237200 1 0 $X=832918 $Y=2231760
X995 2327 2329 2 4 2366 XNOR2X2 $T=933900 2348080 1 0 $X=933898 $Y=2342640
X996 2426 2425 2 4 2445 XNOR2X2 $T=956340 2348080 0 0 $X=956338 $Y=2347678
X997 2439 2440 2 4 2597 XNOR2X2 $T=959640 2368240 0 0 $X=959638 $Y=2367838
X998 2650 2667 2 4 2332 XNOR2X2 $T=1021680 2267440 1 180 $X=1014420 $Y=2267038
X999 2673 2692 2 4 2671 XNOR2X2 $T=1029600 2348080 0 180 $X=1022340 $Y=2342640
X1000 2881 2865 2 4 2807 XNOR2X2 $T=1073820 2317840 0 180 $X=1066560 $Y=2312400
X1001 3037 3026 2 4 2906 XNOR2X2 $T=1113420 2317840 0 180 $X=1106160 $Y=2312400
X1002 3102 3094 2 4 3001 XNOR2X2 $T=1131240 2317840 1 180 $X=1123980 $Y=2317438
X1003 3478 3479 2 4 3497 XNOR2X2 $T=1213080 2277520 0 0 $X=1213078 $Y=2277118
X1004 3930 177 2 4 4065 XNOR2X2 $T=1323300 2287600 0 0 $X=1323298 $Y=2287198
X1005 3985 180 2 4 186 XNOR2X2 $T=1335840 2277520 1 0 $X=1335838 $Y=2272080
X1006 4100 188 2 4 185 XNOR2X2 $T=1364220 2368240 0 180 $X=1356960 $Y=2362800
X1007 6217 6219 2 4 373 XNOR2X2 $T=1910700 2327920 0 0 $X=1910698 $Y=2327518
X1008 6221 6279 2 4 6299 XNOR2X2 $T=1924560 2398480 0 0 $X=1924558 $Y=2398078
X1009 6321 6301 2 4 383 XNOR2X2 $T=1937760 2287600 0 0 $X=1937758 $Y=2287198
X1010 7203 7200 2 4 443 XNOR2X2 $T=2185920 2247280 1 180 $X=2178660 $Y=2246878
X1011 7508 7511 2 4 459 XNOR2X2 $T=2269740 2247280 0 0 $X=2269738 $Y=2246878
X1012 2979 2958 4 2 2957 XOR2X1 $T=1100880 2297680 1 180 $X=1095600 $Y=2297278
X1013 4140 4158 4 2 4163 XOR2X1 $T=1374780 2348080 1 0 $X=1374778 $Y=2342640
X1014 4195 4193 4 2 194 XOR2X1 $T=1387980 2348080 0 180 $X=1382700 $Y=2342640
X1015 4235 4221 4 2 198 XOR2X1 $T=1398540 2388400 1 180 $X=1393260 $Y=2387998
X1016 4291 4281 4 2 203 XOR2X1 $T=1406460 2388400 1 180 $X=1401180 $Y=2387998
X1017 250 4641 4 2 252 XOR2X1 $T=1514040 2237200 1 0 $X=1514038 $Y=2231760
X1018 4706 4705 4 2 4382 XOR2X1 $T=1523940 2287600 1 180 $X=1518660 $Y=2287198
X1019 4792 4791 4 2 4729 XOR2X1 $T=1545060 2247280 1 180 $X=1539780 $Y=2246878
X1020 4802 4764 4 2 4645 XOR2X1 $T=1547700 2267440 1 180 $X=1542420 $Y=2267038
X1021 281 277 4 2 5032 XOR2X1 $T=1613040 2257360 1 180 $X=1607760 $Y=2256958
X1022 273 5157 4 2 5188 XOR2X1 $T=1643400 2247280 1 0 $X=1643398 $Y=2241840
X1023 274 322 4 2 5465 XOR2X1 $T=1716660 2297680 0 0 $X=1716658 $Y=2297278
X1024 271 5482 4 2 5633 XOR2X1 $T=1754280 2368240 1 0 $X=1754278 $Y=2362800
X1025 275 5628 4 2 5649 XOR2X1 $T=1760880 2398480 0 0 $X=1760878 $Y=2398078
X1026 329 5717 4 2 5863 XOR2X1 $T=1785300 2358160 1 0 $X=1785298 $Y=2352720
X1027 5757 5817 4 2 5830 XOR2X1 $T=1801140 2368240 1 0 $X=1801138 $Y=2362800
X1028 348 5924 4 2 6046 XOR2X1 $T=1844040 2378320 1 0 $X=1844038 $Y=2372880
X1029 362 6062 4 2 6074 XOR2X1 $T=1872420 2388400 0 0 $X=1872418 $Y=2387998
X1030 6235 6356 4 2 6443 XOR2X1 $T=1957560 2388400 0 0 $X=1957558 $Y=2387998
X1031 342 6647 4 2 6794 XOR2X1 $T=2028840 2388400 0 0 $X=2028838 $Y=2387998
X1032 6137 6709 4 2 6771 XOR2X1 $T=2052600 2307760 1 0 $X=2052598 $Y=2302320
X1033 434 7012 4 2 6994 XOR2X1 $T=2126520 2408560 0 180 $X=2121240 $Y=2403120
X1034 7283 7282 4 2 450 XOR2X1 $T=2207700 2247280 1 180 $X=2202420 $Y=2246878
X1035 7396 7381 4 2 454 XOR2X1 $T=2245320 2257360 0 180 $X=2240040 $Y=2251920
X1036 7625 7626 4 2 461 XOR2X1 $T=2304060 2247280 0 0 $X=2304058 $Y=2246878
X1037 7817 7794 4 2 464 XOR2X1 $T=2354220 2267440 0 0 $X=2354218 $Y=2267038
X1038 8490 8489 4 2 506 XOR2X1 $T=2531100 2247280 0 0 $X=2531098 $Y=2246878
X1039 1638 2 1660 1724 4 NOR2BX1 $T=755040 2338000 0 180 $X=752400 $Y=2332560
X1040 2653 2 2731 2845 4 NOR2BX1 $T=1063920 2388400 1 0 $X=1063918 $Y=2382960
X1041 2907 2 2908 3002 4 NOR2BX1 $T=1087020 2398480 1 0 $X=1087018 $Y=2393040
X1042 3218 2 3259 3258 4 NOR2BX1 $T=1168200 2307760 0 0 $X=1168198 $Y=2307358
X1043 6142 2 6111 6134 4 NOR2BX1 $T=1895520 2368240 1 180 $X=1892880 $Y=2367838
X1044 29 30 1557 1573 2 4 1576 ADDFX2 $T=700920 2237200 0 0 $X=700918 $Y=2236798
X1045 34 1592 1576 1574 2 4 1559 ADDFX2 $T=724020 2267440 0 180 $X=710160 $Y=2262000
X1046 37 1640 35 1543 2 4 1610 ADDFX2 $T=737880 2237200 1 180 $X=724020 $Y=2236798
X1047 36 38 1655 1672 2 4 1671 ADDFX2 $T=734580 2277520 0 0 $X=734578 $Y=2277118
X1048 1573 1656 1671 1673 2 4 1657 ADDFX2 $T=735240 2277520 1 0 $X=735238 $Y=2272080
X1049 38 42 40 1655 2 4 1592 ADDFX2 $T=749760 2267440 0 180 $X=735900 $Y=2262000
X1050 33 39 41 1683 2 4 1656 ADDFX2 $T=736560 2257360 1 0 $X=736558 $Y=2251920
X1051 42 44 43 1557 2 4 1640 ADDFX2 $T=760980 2237200 1 180 $X=747120 $Y=2236798
X1052 1887 1683 1672 1738 2 4 1736 ADDFX2 $T=770880 2287600 0 180 $X=757020 $Y=2282160
X1053 39 43 1977 1981 2 4 1887 ADDFX2 $T=828300 2277520 0 0 $X=828298 $Y=2277118
X1054 1981 2048 2058 2059 2 4 2076 ADDFX2 $T=846120 2287600 1 0 $X=846118 $Y=2282160
X1055 43 40 2077 2079 2 4 2058 ADDFX2 $T=852720 2277520 1 0 $X=852718 $Y=2272080
X1056 2149 2111 2079 2104 2 4 2089 ADDFX2 $T=882420 2287600 0 180 $X=868560 $Y=2282160
X1057 44 40 38 2147 2 4 2149 ADDFX2 $T=876480 2277520 0 0 $X=876478 $Y=2277118
X1058 42 39 2147 2172 2 4 2168 ADDFX2 $T=905520 2287600 0 180 $X=891660 $Y=2282160
X1059 101 100 98 2674 2 4 2765 ADDFX2 $T=1071180 2247280 0 180 $X=1057320 $Y=2241840
X1060 106 104 102 2866 2 4 2690 ADDFX2 $T=1094280 2247280 1 180 $X=1080420 $Y=2246878
X1061 110 108 105 2918 2 4 2809 ADDFX2 $T=1102200 2237200 0 180 $X=1088340 $Y=2231760
X1062 117 116 113 2937 2 4 2922 ADDFX2 $T=1117380 2247280 0 180 $X=1103520 $Y=2241840
X1063 125 123 122 3126 2 4 3083 ADDFX2 $T=1155660 2237200 1 180 $X=1141800 $Y=2236798
X1064 208 210 4341 213 2 4 4328 ADDFX2 $T=1411740 2287600 1 0 $X=1411738 $Y=2282160
X1065 4395 217 4364 215 2 4 214 ADDFX2 $T=1439460 2307760 0 180 $X=1425600 $Y=2302320
X1066 212 197 218 4378 2 4 4364 ADDFX2 $T=1444740 2277520 1 180 $X=1430880 $Y=2277118
X1067 4378 222 4463 227 2 4 229 ADDFX2 $T=1446720 2327920 0 0 $X=1446718 $Y=2327518
X1068 4473 231 4475 4464 2 4 224 ADDFX2 $T=1466520 2297680 1 180 $X=1452660 $Y=2297278
X1069 197 205 228 4473 2 4 4463 ADDFX2 $T=1467840 2277520 0 180 $X=1453980 $Y=2272080
X1070 205 201 234 4518 2 4 4475 ADDFX2 $T=1459920 2267440 1 0 $X=1459918 $Y=2262000
X1071 4518 242 4550 237 2 4 4462 ADDFX2 $T=1494240 2267440 1 180 $X=1480380 $Y=2267038
X1072 201 195 240 4552 2 4 4550 ADDFX2 $T=1496880 2277520 1 180 $X=1483020 $Y=2277118
X1073 4552 241 4586 245 2 4 246 ADDFX2 $T=1484340 2327920 0 0 $X=1484338 $Y=2327518
X1074 195 209 244 4590 2 4 4586 ADDFX2 $T=1485000 2317840 0 0 $X=1484998 $Y=2317438
X1075 209 211 238 4702 2 4 4689 ADDFX2 $T=1510080 2327920 0 0 $X=1510078 $Y=2327518
X1076 4590 251 4689 4708 2 4 256 ADDFX2 $T=1511400 2338000 0 0 $X=1511398 $Y=2337598
X1077 4881 265 4855 4794 2 4 4824 ADDFX2 $T=1563540 2287600 1 180 $X=1549680 $Y=2287198
X1078 277 274 4903 4882 2 4 4886 ADDFX2 $T=1578060 2277520 0 180 $X=1564200 $Y=2272080
X1079 281 277 270 4888 2 4 4855 ADDFX2 $T=1578060 2307760 0 180 $X=1564200 $Y=2302320
X1080 270 265 271 4889 2 4 4803 ADDFX2 $T=1578060 2368240 0 180 $X=1564200 $Y=2362800
X1081 281 270 273 4902 2 4 4901 ADDFX2 $T=1580700 2247280 0 180 $X=1566840 $Y=2241840
X1082 273 270 274 4904 2 4 4878 ADDFX2 $T=1580700 2317840 1 180 $X=1566840 $Y=2317438
X1083 277 274 265 4780 2 4 4885 ADDFX2 $T=1580700 2358160 0 180 $X=1566840 $Y=2352720
X1084 274 271 275 272 2 4 4883 ADDFX2 $T=1580700 2398480 1 180 $X=1566840 $Y=2398078
X1085 211 210 289 5067 2 4 5063 ADDFX2 $T=1603140 2307760 1 0 $X=1603138 $Y=2302320
X1086 4702 286 5063 5068 2 4 5048 ADDFX2 $T=1603800 2327920 0 0 $X=1603798 $Y=2327518
X1087 210 217 295 5154 2 4 5169 ADDFX2 $T=1634820 2307760 1 0 $X=1634818 $Y=2302320
X1088 5067 5150 5169 5159 2 4 5096 ADDFX2 $T=1634820 2327920 0 0 $X=1634818 $Y=2327518
X1089 5154 296 5187 299 2 4 5170 ADDFX2 $T=1639440 2348080 0 0 $X=1639438 $Y=2347678
X1090 217 222 300 5218 2 4 5187 ADDFX2 $T=1640100 2277520 0 0 $X=1640098 $Y=2277118
X1091 5218 307 5322 5313 2 4 298 ADDFX2 $T=1679040 2287600 0 0 $X=1679038 $Y=2287198
X1092 5351 5345 5326 5323 2 4 5312 ADDFX2 $T=1699500 2327920 1 180 $X=1685640 $Y=2327518
X1093 222 231 313 5351 2 4 5322 ADDFX2 $T=1686300 2277520 0 0 $X=1686298 $Y=2277118
X1094 231 242 314 5359 2 4 5326 ADDFX2 $T=1686960 2307760 1 0 $X=1686958 $Y=2302320
X1095 5442 323 5359 5422 2 4 5406 ADDFX2 $T=1723920 2327920 0 180 $X=1710060 $Y=2322480
X1096 5483 329 5453 5519 2 4 5524 ADDFX2 $T=1727880 2358160 1 0 $X=1727878 $Y=2352720
X1097 5502 316 5535 5546 2 4 5523 ADDFX2 $T=1733160 2327920 1 0 $X=1733158 $Y=2322480
X1098 314 286 5516 5631 2 4 5601 ADDFX2 $T=1753620 2317840 0 0 $X=1753618 $Y=2317438
X1099 6691 403 5280 6730 2 4 6710 ADDFX2 $T=2036760 2277520 1 0 $X=2036758 $Y=2272080
X1100 6736 6662 6771 6787 2 4 6789 ADDFX2 $T=2050620 2297680 0 0 $X=2050618 $Y=2297278
X1101 6137 391 6662 6801 2 4 6865 ADDFX2 $T=2055900 2348080 1 0 $X=2055898 $Y=2342640
X1102 6844 6825 6770 6804 2 4 6802 ADDFX2 $T=2081640 2338000 0 180 $X=2067780 $Y=2332560
X1103 6979 6869 6042 7006 2 4 6855 ADDFX2 $T=2110020 2388400 1 0 $X=2110018 $Y=2382960
X1104 6137 5266 6737 6991 2 4 6979 ADDFX2 $T=2127180 2348080 1 180 $X=2113320 $Y=2347678
X1105 6844 7037 6868 7075 2 4 7068 ADDFX2 $T=2134440 2388400 1 0 $X=2134438 $Y=2382960
X1106 6732 7170 7183 7185 2 4 448 ADDFX2 $T=2172060 2378320 0 0 $X=2172058 $Y=2377918
X1107 7168 6868 7049 7208 2 4 7183 ADDFX2 $T=2176020 2368240 0 0 $X=2176018 $Y=2367838
X1108 6737 7206 7186 7170 2 4 7179 ADDFX2 $T=2190540 2358160 1 180 $X=2176680 $Y=2357758
X1109 5508 7037 7151 7239 2 4 7285 ADDFX2 $T=2186580 2338000 1 0 $X=2186578 $Y=2332560
X1110 5508 5244 7151 7240 2 4 7272 ADDFX2 $T=2187240 2348080 0 0 $X=2187238 $Y=2347678
X1111 6042 7186 7285 7289 2 4 7302 ADDFX2 $T=2197800 2317840 0 0 $X=2197798 $Y=2317438
X1112 6732 7049 7337 7346 2 4 7348 ADDFX2 $T=2214960 2327920 0 0 $X=2214958 $Y=2327518
X1113 7206 7323 7239 7347 2 4 7337 ADDFX2 $T=2215620 2338000 1 0 $X=2215618 $Y=2332560
X1114 7323 5280 5709 7397 2 4 7379 ADDFX2 $T=2232780 2368240 0 0 $X=2232778 $Y=2367838
X1115 7397 7657 7641 7676 2 4 7672 ADDFX2 $T=2308680 2378320 1 0 $X=2308678 $Y=2372880
X1116 7401 7336 7672 7686 2 4 7656 ADDFX2 $T=2309340 2338000 0 0 $X=2309338 $Y=2337598
X1117 5988 7137 5942 7687 2 4 7657 ADDFX2 $T=2309340 2388400 1 0 $X=2309338 $Y=2382960
X1118 7228 5508 7687 7742 2 4 7845 ADDFX2 $T=2331780 2388400 0 0 $X=2331778 $Y=2387998
X1119 5709 7323 6059 7771 2 4 7768 ADDFX2 $T=2333100 2368240 1 0 $X=2333098 $Y=2362800
X1120 7641 7742 7768 7772 2 4 7790 ADDFX2 $T=2335080 2358160 0 0 $X=2335078 $Y=2357758
X1121 7845 7850 6790 7832 2 4 7864 ADDFX2 $T=2362140 2388400 0 0 $X=2362138 $Y=2387998
X1122 5942 5988 6786 8025 2 4 8038 ADDFX2 $T=2401740 2378320 1 0 $X=2401738 $Y=2372880
X1123 8025 7558 8069 8083 2 4 8057 ADDFX2 $T=2419560 2368240 0 0 $X=2419558 $Y=2367838
X1124 7850 7228 8084 8087 2 4 8069 ADDFX2 $T=2422200 2398480 0 0 $X=2422198 $Y=2398078
X1125 6731 5709 6059 8171 2 4 8174 ADDFX2 $T=2440020 2368240 1 0 $X=2440018 $Y=2362800
X1126 6786 5942 7558 8232 2 4 8222 ADDFX2 $T=2459160 2378320 0 0 $X=2459158 $Y=2377918
X1127 8171 8068 8222 8235 2 4 8234 ADDFX2 $T=2461140 2358160 0 0 $X=2461138 $Y=2357758
X1128 8252 8232 8235 8283 2 4 8287 ADDFX2 $T=2477640 2338000 1 0 $X=2477638 $Y=2332560
X1129 472 8297 8285 8313 2 4 8314 ADDFX2 $T=2487540 2317840 1 0 $X=2487538 $Y=2312400
X1130 8084 6732 6772 8285 2 4 8252 ADDFX2 $T=2501400 2348080 0 180 $X=2487540 $Y=2342640
X1131 6786 7850 8068 8378 2 4 8465 ADDFX2 $T=2498100 2378320 1 0 $X=2498098 $Y=2372880
X1132 6772 6790 8378 8546 2 4 8611 ADDFX2 $T=2531760 2348080 1 0 $X=2531758 $Y=2342640
X1133 8418 8308 8465 8556 2 4 8574 ADDFX2 $T=2535060 2358160 0 0 $X=2535058 $Y=2357758
X1134 2766 2756 4 2 2733 XNOR2X1 $T=1048080 2307760 0 180 $X=1042800 $Y=2302320
X1135 3280 3254 4 2 3295 XNOR2X1 $T=1173480 2338000 0 0 $X=1173478 $Y=2337598
X1136 3319 3318 4 2 3308 XNOR2X1 $T=1186680 2317840 1 180 $X=1181400 $Y=2317438
X1137 3574 3582 4 2 3597 XNOR2X1 $T=1236180 2317840 0 0 $X=1236178 $Y=2317438
X1138 3619 3624 4 2 3640 XNOR2X1 $T=1244100 2317840 1 0 $X=1244098 $Y=2312400
X1139 3685 3687 4 2 3744 XNOR2X1 $T=1255980 2297680 1 0 $X=1255978 $Y=2292240
X1140 3682 3708 4 2 3694 XNOR2X1 $T=1265220 2267440 1 180 $X=1259940 $Y=2267038
X1141 4181 4182 4 2 193 XNOR2X1 $T=1386000 2247280 0 180 $X=1380720 $Y=2241840
X1142 4385 4122 4 2 219 XNOR2X1 $T=1434840 2338000 1 0 $X=1434838 $Y=2332560
X1143 4658 248 4 2 4183 XNOR2X1 $T=1511400 2368240 0 180 $X=1506120 $Y=2362800
X1144 5099 5100 4 2 292 XNOR2X1 $T=1623600 2388400 1 0 $X=1623598 $Y=2382960
X1145 5249 5259 4 2 305 XNOR2X1 $T=1667820 2388400 0 0 $X=1667818 $Y=2387998
X1146 340 343 4 2 5833 XNOR2X1 $T=1803780 2388400 0 0 $X=1803778 $Y=2387998
X1147 345 347 4 2 5986 XNOR2X1 $T=1814340 2408560 1 0 $X=1814338 $Y=2403120
X1148 5695 5889 4 2 5910 XNOR2X1 $T=1824900 2327920 0 0 $X=1824898 $Y=2327518
X1149 5908 5912 4 2 5931 XNOR2X1 $T=1830180 2348080 0 0 $X=1830178 $Y=2347678
X1150 335 355 4 2 6034 XNOR2X1 $T=1840740 2348080 0 0 $X=1840738 $Y=2347678
X1151 354 356 4 2 6045 XNOR2X1 $T=1843380 2338000 0 0 $X=1843378 $Y=2337598
X1152 6099 6147 4 2 368 XNOR2X1 $T=1898160 2338000 1 180 $X=1892880 $Y=2337598
X1153 6266 6287 4 2 6304 XNOR2X1 $T=1929180 2358160 0 0 $X=1929178 $Y=2357758
X1154 3959 6427 4 2 395 XNOR2X1 $T=1963500 2237200 1 0 $X=1963498 $Y=2231760
X1155 6949 6946 4 2 6959 XNOR2X1 $T=2102100 2338000 1 0 $X=2102098 $Y=2332560
X1156 7114 7113 4 2 439 XNOR2X1 $T=2154240 2247280 0 0 $X=2154238 $Y=2246878
X1157 7995 8072 4 2 477 XNOR2X1 $T=2428800 2257360 0 0 $X=2428798 $Y=2256958
X1158 8450 8467 4 2 8578 XNOR2X1 $T=2544300 2307760 1 0 $X=2544298 $Y=2302320
X1159 335 5345 4 5345 2 5688 5691 337 OAI221XL $T=1775400 2257360 1 0 $X=1775398 $Y=2251920
X1160 505 8461 4 503 2 8473 8472 8474 OAI221XL $T=2533080 2267440 1 180 $X=2528460 $Y=2267038
X1161 62 1977 44 2 4 2048 ADDHXL $T=836220 2277520 1 0 $X=836218 $Y=2272080
X1162 41 2077 42 2 4 2111 ADDHXL $T=858660 2257360 0 0 $X=858658 $Y=2256958
X1163 38 2296 43 2 4 2350 ADDHXL $T=933240 2317840 1 0 $X=933238 $Y=2312400
X1164 2441 2352 40 2 4 2436 ADDHXL $T=966900 2317840 0 180 $X=959640 $Y=2312400
X1165 204 4278 211 2 4 4318 ADDHXL $T=1413060 2327920 0 0 $X=1413058 $Y=2327518
X1166 204 4341 212 2 4 4395 ADDHXL $T=1417680 2277520 1 0 $X=1417678 $Y=2272080
X1167 241 5442 242 2 4 5453 ADDHXL $T=1712700 2317840 0 0 $X=1712698 $Y=2317438
X1168 251 5483 241 2 4 5535 ADDHXL $T=1731840 2338000 1 0 $X=1731838 $Y=2332560
X1169 286 5502 251 2 4 5516 ADDHXL $T=1743720 2317840 1 180 $X=1736460 $Y=2317438
X1170 6736 6770 6691 2 4 6838 ADDHXL $T=2053260 2338000 0 0 $X=2053258 $Y=2337598
X1171 5244 7037 391 2 4 7089 ADDHXL $T=2129160 2327920 0 0 $X=2129158 $Y=2327518
X1172 2 165 3741 3743 4 NOR2XL $T=1275780 2237200 0 0 $X=1275778 $Y=2236798
X1173 2 170 172 3800 4 NOR2XL $T=1292280 2237200 1 180 $X=1290300 $Y=2236798
X1174 2 195 192 4145 4 NOR2XL $T=1377420 2317840 1 180 $X=1375440 $Y=2317438
X1175 2 339 316 5712 4 NOR2XL $T=1782000 2287600 0 0 $X=1781998 $Y=2287198
X1176 2 5150 329 5737 4 NOR2XL $T=1795200 2317840 1 0 $X=1795198 $Y=2312400
X1177 2 391 5106 6589 4 NOR2XL $T=2010360 2277520 0 180 $X=2008380 $Y=2272080
X1178 2 7719 472 8461 4 NOR2XL $T=2510640 2297680 1 0 $X=2510638 $Y=2292240
X1179 2 7719 8424 501 4 NOR2XL $T=2521200 2287600 0 0 $X=2521198 $Y=2287198
X1180 2 8473 502 8449 4 NOR2XL $T=2523840 2257360 0 0 $X=2523838 $Y=2256958
X1181 3843 172 170 4 2 3794 XOR3X2 $T=1298880 2267440 1 180 $X=1287000 $Y=2267038
X1182 5428 5422 5524 4 2 334 XOR3X2 $T=1735140 2408560 1 0 $X=1735138 $Y=2403120
X1183 5266 403 6589 4 2 402 XOR3X2 $T=2014980 2257360 1 180 $X=2003100 $Y=2256958
X1184 6662 6648 6621 4 2 405 XOR3X2 $T=2028180 2307760 0 180 $X=2016300 $Y=2302320
X1185 6789 6730 6761 4 2 414 XOR3X2 $T=2064480 2257360 0 180 $X=2052600 $Y=2251920
X1186 3720 3684 2 3675 4 160 AOI21XL $T=1257300 2378320 0 180 $X=1254660 $Y=2372880
X1187 3751 3691 2 3747 4 3718 AOI21XL $T=1275780 2247280 1 180 $X=1273140 $Y=2246878
X1188 3691 3743 2 3763 4 3810 AOI21XL $T=1275780 2247280 1 0 $X=1275778 $Y=2241840
X1189 6134 370 2 6218 4 6232 AOI21XL $T=1910040 2378320 1 0 $X=1910038 $Y=2372880
X1190 370 6222 2 6252 4 6282 AOI21XL $T=1920600 2408560 0 0 $X=1920598 $Y=2408158
X1191 370 6269 2 6277 4 6286 AOI21XL $T=1924560 2368240 0 0 $X=1924558 $Y=2367838
X1192 6267 370 2 6263 4 6398 AOI21XL $T=1952940 2368240 0 0 $X=1952938 $Y=2367838
X1193 8449 493 2 8474 4 8489 AOI21XL $T=2529780 2257360 1 0 $X=2529778 $Y=2251920
X1194 1900 56 1898 4 1885 2 OAI2BB1X1 $T=811140 2257360 0 0 $X=811138 $Y=2256958
X1195 3475 3595 3581 4 3582 2 OAI2BB1X1 $T=1240800 2297680 1 180 $X=1237500 $Y=2297278
X1196 3961 180 3897 4 3976 2 OAI2BB1X1 $T=1331220 2317840 1 0 $X=1331218 $Y=2312400
X1197 4229 200 4208 4 4181 2 OAI2BB1X1 $T=1392600 2237200 1 180 $X=1389300 $Y=2236798
X1198 5278 5283 5294 4 5314 2 OAI2BB1X1 $T=1675740 2398480 1 0 $X=1675738 $Y=2393040
X1199 335 5345 5647 4 5606 2 OAI2BB1X1 $T=1768140 2267440 0 0 $X=1768138 $Y=2267038
X1200 319 5651 5658 4 5677 2 OAI2BB1X1 $T=1770120 2378320 0 0 $X=1770118 $Y=2377918
X1201 6253 376 6232 4 6147 2 OAI2BB1X1 $T=1920600 2378320 0 180 $X=1917300 $Y=2372880
X1202 6303 376 6282 4 6279 2 OAI2BB1X1 $T=1931160 2408560 1 180 $X=1927860 $Y=2408158
X1203 6602 6589 6619 4 6621 2 OAI2BB1X1 $T=2009040 2277520 0 0 $X=2009038 $Y=2277118
X1204 2108 4 2107 2 2090 NAND2BXL $T=873180 2358160 0 180 $X=870540 $Y=2352720
X1205 2676 4 2672 2 2673 NAND2BXL $T=1024320 2307760 0 180 $X=1021680 $Y=2302320
X1206 2919 4 2920 2 2881 NAND2BXL $T=1084380 2297680 1 180 $X=1081740 $Y=2297278
X1207 3003 4 2997 2 2979 NAND2BXL $T=1102860 2267440 1 180 $X=1100220 $Y=2267038
X1208 3091 4 3081 2 3037 NAND2BXL $T=1126620 2267440 0 180 $X=1123980 $Y=2262000
X1209 2999 4 2959 2 3100 NAND2BXL $T=1126620 2398480 1 0 $X=1126618 $Y=2393040
X1210 3197 4 3204 2 3202 NAND2BXL $T=1153680 2277520 0 180 $X=1151040 $Y=2272080
X1211 3259 4 3310 2 3280 NAND2BXL $T=1189320 2307760 1 0 $X=1189318 $Y=2302320
X1212 3334 4 3336 2 3319 NAND2BXL $T=1189980 2287600 1 0 $X=1189978 $Y=2282160
X1213 3477 4 3471 2 3450 NAND2BXL $T=1213080 2277520 0 180 $X=1210440 $Y=2272080
X1214 155 4 153 2 3574 NAND2BXL $T=1238820 2247280 0 180 $X=1236180 $Y=2241840
X1215 3880 4 3881 2 3930 NAND2BXL $T=1301520 2287600 1 0 $X=1301518 $Y=2282160
X1216 4737 4 4714 2 4676 NAND2BXL $T=1526580 2317840 1 180 $X=1523940 $Y=2317438
X1217 4877 4 4880 2 269 NAND2BXL $T=1570800 2237200 0 180 $X=1568160 $Y=2231760
X1218 5062 4 5046 2 287 NAND2BXL $T=1610400 2388400 0 180 $X=1607760 $Y=2382960
X1219 5082 4 5098 2 5099 NAND2BXL $T=1623600 2378320 0 180 $X=1620960 $Y=2372880
X1220 231 4 311 2 5424 NAND2BXL $T=1691580 2267440 0 0 $X=1691578 $Y=2267038
X1221 5405 4 5404 2 317 NAND2BXL $T=1708740 2378320 0 180 $X=1706100 $Y=2372880
X1222 5607 4 5708 2 5630 NAND2BXL $T=1783320 2348080 1 180 $X=1780680 $Y=2347678
X1223 5150 4 338 2 5740 NAND2BXL $T=1789260 2267440 0 0 $X=1789258 $Y=2267038
X1224 5607 4 5676 2 5832 NAND2BXL $T=1810380 2358160 0 0 $X=1810378 $Y=2357758
X1225 6081 4 6028 2 6099 NAND2BXL $T=1879680 2348080 0 0 $X=1879678 $Y=2347678
X1226 5993 4 6015 2 6221 NAND2BXL $T=1895520 2398480 0 0 $X=1895518 $Y=2398078
X1227 6461 6464 4 2 CLKBUFX3 $T=1971420 2297680 0 0 $X=1971418 $Y=2297278
X1228 3800 3810 170 172 2 4 3825 AOI2BB2X1 $T=1288980 2247280 1 0 $X=1288978 $Y=2241840
X1229 260 4780 4803 4767 2 4 4781 ADDFHX1 $T=1533840 2358160 0 0 $X=1533838 $Y=2357758
X1230 278 4889 4883 268 2 4 4769 ADDFHX1 $T=1576740 2388400 1 180 $X=1561560 $Y=2387998
X1231 5106 6736 6844 6869 2 4 6847 ADDFHX1 $T=2075700 2378320 1 0 $X=2075698 $Y=2372880
X1232 6801 6847 6868 6853 2 4 6866 ADDFHX1 $T=2076360 2388400 0 0 $X=2076358 $Y=2387998
X1233 6838 6865 6737 6867 2 4 6870 ADDFHX1 $T=2080980 2348080 0 0 $X=2080978 $Y=2347678
X1234 6991 7049 7068 7071 2 4 7011 ADDFHX1 $T=2129160 2398480 1 0 $X=2129158 $Y=2393040
X1235 5988 7168 7186 7363 2 4 7364 ADDFHX1 $T=2217600 2388400 0 0 $X=2217598 $Y=2387998
X1236 5314 4 5340 2 5341 5346 NAND3X1 $T=1692900 2398480 1 0 $X=1692898 $Y=2393040
X1237 7181 4 7182 2 7184 444 NAND3X1 $T=2179320 2408560 1 0 $X=2179318 $Y=2403120
X1238 7476 4 7478 2 7479 7480 NAND3X1 $T=2260500 2368240 1 0 $X=2260498 $Y=2362800
X1239 8173 4 8170 2 8101 8186 NAND3X1 $T=2455200 2338000 0 0 $X=2455198 $Y=2337598
X1240 6731 6732 6059 8308 4 2 8297 CMPR32X1 $T=2484900 2358160 0 0 $X=2484898 $Y=2357758
X1241 4101 4102 4009 4 4070 2 AOI2BB1X2 $T=1364220 2378320 0 180 $X=1359600 $Y=2372880
X1242 271 4888 4878 4854 2 4 4789 ADDFHX2 $T=1581360 2317840 0 180 $X=1558920 $Y=2312400
X1243 275 4904 4885 4777 2 4 4851 ADDFHX2 $T=1584000 2338000 0 180 $X=1561560 $Y=2332560
X1244 5266 7137 7150 7151 2 4 7168 ADDFHX2 $T=2148300 2338000 0 0 $X=2148298 $Y=2337598
X1245 5106 5280 7089 7150 2 4 7206 ADDFHX2 $T=2150280 2327920 0 0 $X=2150278 $Y=2327518
X1246 7208 7302 7316 7305 2 4 7167 ADDFHX2 $T=2197140 2287600 0 0 $X=2197138 $Y=2287198
X1247 7289 7336 7348 7352 2 4 7315 ADDFHX2 $T=2210340 2307760 1 0 $X=2210338 $Y=2302320
X1248 7240 7379 7316 7401 2 4 7451 ADDFHX2 $T=2225520 2358160 1 0 $X=2225518 $Y=2352720
X1249 7347 7364 7316 7403 2 4 7410 ADDFHX2 $T=2226180 2317840 0 0 $X=2226178 $Y=2317438
X1250 7346 7410 6790 7464 2 4 7450 ADDFHX2 $T=2236080 2297680 0 0 $X=2236078 $Y=2297278
X1251 7228 7272 7363 7477 2 4 7510 ADDFHX2 $T=2247960 2398480 1 0 $X=2247958 $Y=2393040
X1252 7336 7403 7571 7574 2 4 7512 ADDFHX2 $T=2272380 2317840 0 0 $X=2272378 $Y=2317438
X1253 6976 7624 7640 7642 2 4 7639 ADDFHX2 $T=2288220 2348080 1 0 $X=2288218 $Y=2342640
X1254 6732 7510 7641 7624 2 4 7571 ADDFHX2 $T=2288220 2368240 1 0 $X=2288218 $Y=2362800
X1255 7719 7480 7656 7654 2 4 7651 ADDFHX2 $T=2332440 2327920 0 180 $X=2310000 $Y=2322480
X1256 6976 7676 7864 7867 2 4 7866 ADDFHX2 $T=2351580 2388400 1 0 $X=2351578 $Y=2382960
X1257 7686 7849 7866 7847 2 4 7818 ADDFHX2 $T=2352240 2327920 0 0 $X=2352238 $Y=2327518
X1258 7832 7882 7867 7896 2 4 7846 ADDFHX2 $T=2359500 2348080 0 0 $X=2359498 $Y=2347678
X1259 7558 6772 7790 7897 2 4 7882 ADDFHX2 $T=2360820 2358160 0 0 $X=2360818 $Y=2357758
X1260 7772 472 7719 8008 2 4 7996 ADDFHX2 $T=2385900 2307760 1 0 $X=2385898 $Y=2302320
X1261 8040 7897 7996 7995 2 4 7946 ADDFHX2 $T=2419560 2297680 0 180 $X=2397120 $Y=2292240
X1262 7771 6976 8038 8041 2 4 8040 ADDFHX2 $T=2398440 2358160 1 0 $X=2398438 $Y=2352720
X1263 7719 8041 7849 8082 2 4 8108 ADDFHX2 $T=2417580 2327920 0 0 $X=2417578 $Y=2327518
X1264 8174 8087 472 8100 2 4 8086 ADDFHX2 $T=2457180 2388400 1 180 $X=2434740 $Y=2387998
X1265 7849 8100 8234 8236 2 4 8215 ADDFHX2 $T=2453220 2327920 1 0 $X=2453218 $Y=2322480
X1266 8057 8008 8108 8123 8072 4 2 ADDFHX4 $T=2422860 2307760 1 0 $X=2422858 $Y=2302320
X1267 94 2 2667 4 CLKINVX3 $T=1024980 2277520 1 0 $X=1024978 $Y=2272080
X1268 4101 2 188 4 CLKINVX3 $T=1364220 2358160 1 180 $X=1362240 $Y=2357758
X1269 197 2 192 4 CLKINVX3 $T=1390620 2277520 1 180 $X=1388640 $Y=2277118
X1270 4363 2 4362 4 CLKINVX3 $T=1429560 2368240 0 180 $X=1427580 $Y=2362800
X1271 209 2 218 4 CLKINVX3 $T=1437480 2247280 1 0 $X=1437478 $Y=2241840
X1272 4412 2 4461 4 CLKINVX3 $T=1453980 2378320 0 0 $X=1453978 $Y=2377918
X1273 244 2 222 4 CLKINVX3 $T=1527240 2267440 1 0 $X=1527238 $Y=2262000
X1274 290 2 5264 4 CLKINVX3 $T=1676400 2388400 1 0 $X=1676398 $Y=2382960
X1275 278 2 319 4 CLKINVX3 $T=1698180 2368240 0 0 $X=1698178 $Y=2367838
X1276 5482 2 5557 4 CLKINVX3 $T=1747680 2297680 1 0 $X=1747678 $Y=2292240
X1277 6002 2 6040 4 CLKINVX3 $T=1853280 2277520 1 180 $X=1851300 $Y=2277118
X1278 5559 2 6137 4 CLKINVX3 $T=1892880 2307760 1 0 $X=1892878 $Y=2302320
X1279 6046 2 6732 4 CLKINVX3 $T=2049960 2378320 0 180 $X=2047980 $Y=2372880
X1280 6794 2 6976 4 CLKINVX3 $T=2099460 2388400 1 0 $X=2099458 $Y=2382960
X1281 7009 2 7053 4 CLKINVX3 $T=2123220 2257360 1 0 $X=2123218 $Y=2251920
X1282 5508 2 6844 4 CLKINVX3 $T=2124540 2368240 0 0 $X=2124538 $Y=2367838
X1283 6137 2 7137 4 CLKINVX3 $T=2133780 2348080 0 0 $X=2133778 $Y=2347678
X1284 5709 2 7049 4 CLKINVX3 $T=2154240 2378320 1 0 $X=2154238 $Y=2372880
X1285 7086 2 442 4 CLKINVX3 $T=2164800 2237200 1 0 $X=2164798 $Y=2231760
X1286 6737 2 7323 4 CLKINVX3 $T=2199120 2368240 1 0 $X=2199118 $Y=2362800
X1287 5942 2 7186 4 CLKINVX3 $T=2218260 2368240 0 0 $X=2218258 $Y=2367838
X1288 7319 2 7381 4 CLKINVX3 $T=2230800 2257360 1 0 $X=2230798 $Y=2251920
X1289 7623 2 7671 4 CLKINVX3 $T=2300760 2277520 1 180 $X=2298780 $Y=2277118
X1290 6732 2 7850 4 CLKINVX3 $T=2385240 2378320 1 0 $X=2385238 $Y=2372880
X1291 6976 2 8068 4 CLKINVX3 $T=2426820 2358160 0 0 $X=2426818 $Y=2357758
X1292 6790 2 8084 4 CLKINVX3 $T=2429460 2408560 1 0 $X=2429458 $Y=2403120
X1293 6731 2 7641 4 CLKINVX3 $T=2486880 2368240 0 0 $X=2486878 $Y=2367838
X1294 7558 2 8418 4 CLKINVX3 $T=2505360 2388400 1 0 $X=2505358 $Y=2382960
X1295 3929 3898 2 4 3946 AND2X1 $T=1322640 2267440 1 0 $X=1322638 $Y=2262000
X1296 4776 4852 2 4 4792 AND2X1 $T=1552980 2257360 0 180 $X=1550340 $Y=2251920
X1297 5219 5151 2 4 5229 AND2X1 $T=1654620 2398480 0 0 $X=1654618 $Y=2398078
X1298 375 6222 2 4 6303 AND2X1 $T=1938420 2408560 1 180 $X=1935780 $Y=2408158
X1299 6284 6191 6234 2 6289 4 AOI2BB1X4 $T=1927200 2317840 0 0 $X=1927198 $Y=2317438
X1300 3596 3594 2 152 154 3581 4 AOI22X1 $T=1240800 2277520 0 180 $X=1237500 $Y=2272080
X1301 5159 5170 2 293 5151 5171 4 AOI22X1 $T=1642740 2398480 1 0 $X=1642738 $Y=2393040
X1302 8475 8516 2 8467 8450 8523 4 AOI22X1 $T=2537040 2307760 1 0 $X=2537038 $Y=2302320
X1303 6710 6694 6713 6692 4 2 6761 OAI2BB2X1 $T=2042700 2267440 1 0 $X=2042698 $Y=2262000
X1304 8068 6731 8418 8424 4 2 8450 ADDFXL $T=2508660 2358160 0 0 $X=2508658 $Y=2357758
X1305 8084 7641 472 8467 4 2 8549 ADDFXL $T=2516580 2327920 1 0 $X=2516578 $Y=2322480
X1306 175 3882 4 2 3898 XNOR2XL $T=1304160 2237200 1 0 $X=1304158 $Y=2231760
X1307 5345 5629 4 2 5645 XNOR2XL $T=1762200 2348080 0 0 $X=1762198 $Y=2347678
X1308 2633 2613 2651 2 4 OR2X4 $T=1014420 2398480 1 0 $X=1014418 $Y=2393040
X1309 2328 182 4066 2 4 OR2X4 $T=1349700 2307760 1 0 $X=1349698 $Y=2302320
X1310 2455 187 4086 2 4 OR2X4 $T=1357620 2297680 0 0 $X=1357618 $Y=2297278
X1311 3239 216 4379 2 4 OR2X4 $T=1430880 2388400 1 0 $X=1430878 $Y=2382960
X1312 2735 220 4409 2 4 OR2X4 $T=1440780 2398480 0 0 $X=1440778 $Y=2398078
X1313 274 322 5444 2 4 OR2X4 $T=1715340 2297680 1 0 $X=1715338 $Y=2292240
X1314 265 5444 5482 2 4 OR2X4 $T=1725900 2297680 1 0 $X=1725898 $Y=2292240
X1315 5507 311 5924 2 4 OR2X4 $T=1836120 2378320 0 0 $X=1836118 $Y=2377918
X1316 3150 358 5990 2 4 OR2X4 $T=1850640 2307760 1 0 $X=1850638 $Y=2302320
X1317 3256 360 6044 2 4 OR2X4 $T=1867140 2327920 0 0 $X=1867138 $Y=2327518
X1318 3159 369 6189 2 4 OR2X4 $T=1898820 2307760 0 0 $X=1898818 $Y=2307358
X1319 3331 377 6260 2 4 OR2X4 $T=1931160 2338000 0 180 $X=1927200 $Y=2332560
X1320 3931 6443 6444 2 4 OR2X4 $T=1968120 2358160 0 0 $X=1968118 $Y=2357758
X1321 336 6678 410 2 4 OR2X4 $T=2037420 2408560 1 0 $X=2037418 $Y=2403120
X1322 7315 7305 7284 2 4 OR2X4 $T=2216280 2277520 1 180 $X=2212320 $Y=2277118
X1323 410 460 7558 2 4 OR2X4 $T=2285580 2408560 1 0 $X=2285578 $Y=2403120
X1324 7639 7574 7643 2 4 OR2X4 $T=2306700 2297680 1 0 $X=2306698 $Y=2292240
X1325 7651 7642 7677 2 4 OR2X4 $T=2325180 2297680 0 0 $X=2325178 $Y=2297278
X1326 469 468 467 2 4 OR2X4 $T=2376000 2237200 0 180 $X=2372040 $Y=2231760
X1327 303 5231 5263 4 2 5280 OAI2BB1X4 $T=1669140 2267440 1 0 $X=1669138 $Y=2262000
X1328 56 1687 4 2 INVX8 $T=801240 2307760 0 180 $X=797280 $Y=2302320
X1329 2612 2616 4 2 INVX8 $T=1005840 2368240 1 180 $X=1001880 $Y=2367838
X1330 6041 6262 4 2 INVX8 $T=1925880 2287600 1 180 $X=1921920 $Y=2287198
X1331 416 6790 4 2 INVX8 $T=2065140 2408560 1 180 $X=2061180 $Y=2408158
X1332 6042 7228 4 2 INVX8 $T=2209680 2398480 0 0 $X=2209678 $Y=2398078
X1333 4119 4117 4067 191 2 4 MX2X4 $T=1365540 2287600 1 0 $X=1365538 $Y=2282160
X1334 6693 336 6678 6772 2 4 MX2X4 $T=2038080 2398480 0 0 $X=2038078 $Y=2398078
X1335 7995 8072 8009 4 8088 8089 2 OAI2BB2X4 $T=2426820 2267440 0 0 $X=2426818 $Y=2267038
X1336 99 111 3024 4 2 NAND2BX2 $T=1108800 2398480 0 0 $X=1108798 $Y=2398078
X1337 5217 5168 5906 4 2 NAND2BX2 $T=1833480 2267440 1 0 $X=1833478 $Y=2262000
X1338 6442 6409 401 4 2 NAND2BX2 $T=1997820 2247280 0 0 $X=1997818 $Y=2246878
X1339 2878 2756 2842 2865 2 4 OAI2BB1X2 $T=1071180 2307760 0 180 $X=1066560 $Y=2302320
X1340 3035 3107 2959 3127 2 4 OAI2BB1X2 $T=1129260 2408560 1 0 $X=1129258 $Y=2403120
X1341 4122 4379 4363 4420 2 4 OAI2BB1X2 $T=1432860 2358160 0 0 $X=1432858 $Y=2357758
X1342 5159 5170 5219 4 2 301 AND3X2 $T=1654620 2408560 1 0 $X=1654618 $Y=2403120
X1343 4234 4215 4 2 4180 XOR2XL $T=1398540 2307760 1 180 $X=1393260 $Y=2307358
X1344 205 204 4 2 4292 XOR2XL $T=1411740 2277520 1 180 $X=1406460 $Y=2277118
X1345 391 5106 4 2 393 XOR2XL $T=1974060 2267440 1 0 $X=1974058 $Y=2262000
X1346 39 2 2441 4 BUFX3 $T=962280 2297680 1 0 $X=962278 $Y=2292240
X1347 2756 2 3019 4 BUFX3 $T=1097580 2297680 1 0 $X=1097578 $Y=2292240
X1348 2616 2 132 4 BUFX3 $T=1178100 2408560 0 0 $X=1178098 $Y=2408158
X1349 3970 2 3959 4 BUFX3 $T=1330560 2257360 1 180 $X=1327920 $Y=2256958
X1350 5188 2 5266 4 BUFX3 $T=1667820 2247280 1 0 $X=1667818 $Y=2241840
X1351 5465 2 5559 4 BUFX3 $T=1721940 2297680 0 0 $X=1721938 $Y=2297278
X1352 7829 2 7819 4 BUFX3 $T=2358180 2307760 1 0 $X=2358178 $Y=2302320
X1353 2189 2151 2196 2 2106 4 2240 2260 AOI221X1 $T=904860 2327920 0 0 $X=904858 $Y=2327518
X1354 5713 5716 5689 2 5708 4 5719 5594 AOI221X1 $T=1783320 2338000 1 0 $X=1783318 $Y=2332560
X1355 303 270 2 4 CLKINVX4 $T=1660560 2247280 1 180 $X=1657920 $Y=2246878
X1356 6461 392 2 4 CLKINVX4 $T=1975380 2297680 0 180 $X=1972740 $Y=2292240
X1357 4220 2 4213 4195 4 NOR2BXL $T=1401180 2327920 1 180 $X=1398540 $Y=2327518
X1358 204 2 205 4234 4 NOR2BXL $T=1401180 2297680 0 0 $X=1401178 $Y=2297278
X1359 231 2 311 5423 4 NOR2BXL $T=1691580 2247280 0 0 $X=1691578 $Y=2246878
X1360 5504 2 5500 332 4 NOR2BXL $T=1741080 2388400 0 0 $X=1741078 $Y=2387998
X1361 5150 2 338 5710 4 NOR2BXL $T=1780020 2267440 0 0 $X=1780018 $Y=2267038
X1362 8122 2 8187 8216 4 NOR2BXL $T=2468400 2257360 0 180 $X=2465760 $Y=2251920
X1363 1643 1622 4 2 1608 1611 AOI2BB1X1 $T=727320 2327920 0 180 $X=724020 $Y=2322480
X1364 5265 5443 4 2 5439 5427 AOI2BB1X1 $T=1717980 2398480 1 180 $X=1714680 $Y=2398078
X1365 335 5688 4 2 5673 5691 AOI2BB1X1 $T=1785960 2257360 0 180 $X=1782660 $Y=2251920
X1366 6821 6863 4 2 6877 6884 AOI2BB1X1 $T=2090220 2297680 1 0 $X=2090218 $Y=2292240
X1367 5648 260 5714 341 4 2 MXI2X1 $T=1780680 2398480 1 0 $X=1780678 $Y=2393040
X1368 313 331 4 330 2 5498 5501 OAI211X1 $T=1735140 2237200 1 180 $X=1731180 $Y=2236798
X1369 2714 2690 2674 4 2 2615 XNOR3X2 $T=1033560 2327920 1 180 $X=1021680 $Y=2327518
X1370 6710 6694 6692 4 2 409 XNOR3X2 $T=2047320 2257360 1 180 $X=2035440 $Y=2256958
X1371 6802 6787 6821 4 2 420 XNOR3X2 $T=2071080 2297680 1 0 $X=2071078 $Y=2292240
X1372 6962 6855 6853 4 2 6947 XNOR3X2 $T=2112000 2398480 0 180 $X=2100120 $Y=2393040
X1373 426 6947 6980 4 2 433 XNOR3X2 $T=2113320 2287600 1 0 $X=2113318 $Y=2282160
X1374 7075 7228 7179 4 2 7138 XNOR3X2 $T=2201100 2398480 1 180 $X=2189220 $Y=2398078
X1375 2960 2 3020 115 114 3011 4 AOI22XL $T=1109460 2277520 0 0 $X=1109458 $Y=2277118
X1376 5829 2 5847 329 5150 5828 4 AOI22XL $T=1808400 2338000 0 180 $X=1805100 $Y=2332560
X1377 5649 5988 4 2 BUFX4 $T=1840740 2398480 0 0 $X=1840738 $Y=2398078
X1378 493 495 4 2 BUFX4 $T=2505360 2237200 1 0 $X=2505358 $Y=2231760
X1379 5423 242 4 5423 320 5438 2 OAI22XL $T=1710720 2247280 0 0 $X=1710718 $Y=2246878
X1380 5470 251 4 5470 326 5498 2 OAI22XL $T=1723260 2247280 1 0 $X=1723258 $Y=2241840
X1381 5710 339 4 5710 340 5650 2 OAI22XL $T=1781340 2277520 0 0 $X=1781338 $Y=2277118
X1382 306 5443 290 4 5427 2 5428 OAI31X1 $T=1718640 2408560 1 180 $X=1714680 $Y=2408158
X1383 5424 242 320 4 5424 2 320 242 5425 OAI222XL $T=1713360 2267440 0 0 $X=1713358 $Y=2267038
X1384 5425 295 321 4 5425 2 295 321 5452 OAI222XL $T=1714680 2267440 1 0 $X=1714678 $Y=2262000
X1385 5452 251 251 4 326 2 5452 326 5522 OAI222XL $T=1722600 2257360 1 0 $X=1722598 $Y=2251920
X1386 5522 313 331 4 5522 2 313 331 5593 OAI222XL $T=1739760 2257360 1 0 $X=1739758 $Y=2251920
X1387 5740 339 5740 4 340 2 340 339 5734 OAI222XL $T=1791900 2267440 0 180 $X=1786620 $Y=2262000
X1388 329 5734 336 4 5734 2 329 336 5688 OAI222XL $T=1787940 2257360 1 0 $X=1787938 $Y=2251920
X1389 5557 333 4 2 5506 AND2X4 $T=1747680 2287600 1 0 $X=1747678 $Y=2282160
X1390 5517 4 5506 5488 2 5507 NAND3X4 $T=1737780 2287600 0 180 $X=1731180 $Y=2282160
X1391 6409 6431 4 387 6440 6449 2 6427 OAI221X2 $T=1964820 2247280 1 0 $X=1964818 $Y=2241840
X1392 5877 349 320 326 2 4 5897 NAND4X4 $T=1831500 2378320 0 180 $X=1820280 $Y=2372880
X1393 4903 273 279 2 4 4881 CMPR22X1 $T=1579380 2287600 1 180 $X=1571460 $Y=2287198
X1394 6648 6709 6691 2 4 6694 CMPR22X1 $T=2046660 2307760 0 180 $X=2038740 $Y=2302320
X1395 94 2668 92 4 93 2687 2 AOI2BB2X4 $T=1022340 2247280 1 0 $X=1022338 $Y=2241840
X1396 7451 7477 6790 7640 4 2 XOR3X4 $T=2254560 2348080 0 0 $X=2254558 $Y=2347678
X1397 8086 8082 8083 8172 4 2 XOR3X4 $T=2432100 2348080 1 0 $X=2432098 $Y=2342640
.ENDS
***************************************
.SUBCKT ICV_56 2 4 41 42 43 44 45 46 47 50 52 54 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 71 72 73 74 75 76 77 78 79 80 81 82 83 84
+ 85 86 87 88 89 90 91 93 94 95 97 98 99 102 103 106 107 108 111 112
+ 114 115 116 117 119 120 123 124 126 127 128 129 130 131 132 134 136 137 138 139
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 195 196 197 198 199 200 201
+ 202 203 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 1248
+ 1249
** N=24561 EP=161 IP=3461 FDC=0
X0 3122 2 2840 4 3120 NAND2X1 $T=1213080 2418640 0 180 $X=1211100 $Y=2413200
X1 60 2 3222 4 3141 NAND2X1 $T=1246740 2418640 1 180 $X=1244760 $Y=2418238
X2 62 2 63 4 3222 NAND2X1 $T=1257300 2418640 0 0 $X=1257298 $Y=2418238
X3 3623 2 3613 4 3588 NAND2X1 $T=1364220 2519440 1 180 $X=1362240 $Y=2519038
X4 3613 2 3624 4 3606 NAND2X1 $T=1364880 2519440 1 0 $X=1364878 $Y=2514000
X5 3626 2 80 4 3605 NAND2X1 $T=1366860 2479120 0 180 $X=1364880 $Y=2473680
X6 3698 2 3623 4 3660 NAND2X1 $T=1379400 2519440 0 180 $X=1377420 $Y=2514000
X7 80 2 3626 4 3657 NAND2X1 $T=1380720 2479120 0 0 $X=1380718 $Y=2478718
X8 3680 2 81 4 3540 NAND2X1 $T=1383360 2428720 0 0 $X=1383358 $Y=2428318
X9 3690 2 3696 4 3631 NAND2X1 $T=1387980 2499280 0 0 $X=1387978 $Y=2498878
X10 82 2 3712 4 3593 NAND2X1 $T=1393920 2438800 1 0 $X=1393918 $Y=2433360
X11 3803 2 3773 4 3624 NAND2X1 $T=1413060 2529520 1 0 $X=1413058 $Y=2524080
X12 85 2 84 4 3770 NAND2X1 $T=1420980 2448880 0 180 $X=1419000 $Y=2443440
X13 86 2 87 4 3874 NAND2X1 $T=1430220 2418640 1 0 $X=1430218 $Y=2413200
X14 3876 2 3878 4 3862 NAND2X1 $T=1431540 2529520 0 0 $X=1431538 $Y=2529118
X15 3878 2 3899 4 3902 NAND2X1 $T=1438140 2529520 1 0 $X=1438138 $Y=2524080
X16 90 2 3904 4 3876 NAND2X1 $T=1442100 2539600 1 180 $X=1440120 $Y=2539198
X17 95 2 93 4 3934 NAND2X1 $T=1455960 2428720 1 180 $X=1453980 $Y=2428318
X18 3995 2 3974 4 3772 NAND2X1 $T=1459260 2519440 1 0 $X=1459258 $Y=2514000
X19 3989 2 4015 4 4032 NAND2X1 $T=1467180 2489200 1 0 $X=1467178 $Y=2483760
X20 4065 2 4015 4 4030 NAND2X1 $T=1469820 2479120 0 180 $X=1467840 $Y=2473680
X21 4033 2 4043 4 3971 NAND2X1 $T=1470480 2559760 1 0 $X=1470478 $Y=2554320
X22 103 2 102 4 4109 NAND2X1 $T=1490280 2448880 1 0 $X=1490278 $Y=2443440
X23 4117 2 4012 4 4120 NAND2X1 $T=1492920 2539600 0 0 $X=1492918 $Y=2539198
X24 106 2 107 4 4170 NAND2X1 $T=1500840 2458960 0 0 $X=1500838 $Y=2458558
X25 4190 2 4185 4 4051 NAND2X1 $T=1509420 2539600 0 0 $X=1509418 $Y=2539198
X26 119 2 4312 4 4192 NAND2X1 $T=1548360 2428720 1 0 $X=1548358 $Y=2423280
X27 120 2 4318 4 4203 NAND2X1 $T=1550340 2549680 0 0 $X=1550338 $Y=2549278
X28 4343 2 4319 4 4220 NAND2X1 $T=1552320 2438800 1 180 $X=1550340 $Y=2438398
X29 4395 2 4361 4 4296 NAND2X1 $T=1568820 2479120 0 0 $X=1568818 $Y=2478718
X30 4407 2 4377 4 4406 NAND2X1 $T=1570800 2539600 0 180 $X=1568820 $Y=2534160
X31 4412 2 4420 4 4403 NAND2X1 $T=1576740 2489200 1 0 $X=1576738 $Y=2483760
X32 4446 2 4407 4 4270 NAND2X1 $T=1580040 2529520 0 180 $X=1578060 $Y=2524080
X33 4377 2 4473 4 136 NAND2X1 $T=1589940 2549680 1 0 $X=1589938 $Y=2544240
X34 4497 2 4488 4 4446 NAND2X1 $T=1594560 2519440 0 180 $X=1592580 $Y=2514000
X35 4559 2 4568 4 4475 NAND2X1 $T=1615680 2529520 1 0 $X=1615678 $Y=2524080
X36 155 2 151 4 152 NAND2X1 $T=1638780 2418640 0 180 $X=1636800 $Y=2413200
X37 4708 2 4646 4 4547 NAND2X1 $T=1649340 2569840 0 180 $X=1647360 $Y=2564400
X38 4739 2 4704 4 4725 NAND2X1 $T=1665840 2549680 0 0 $X=1665838 $Y=2549278
X39 4774 2 4792 4 4678 NAND2X1 $T=1679700 2549680 1 0 $X=1679698 $Y=2544240
X40 4890 2 4840 4 4795 NAND2X1 $T=1700160 2559760 1 180 $X=1698180 $Y=2559358
X41 5072 2 4954 4 5088 NAND2X1 $T=1766160 2529520 1 0 $X=1766158 $Y=2524080
X42 5102 2 177 4 5128 NAND2X1 $T=1770120 2438800 1 0 $X=1770118 $Y=2433360
X43 5157 2 178 4 5233 NAND2X1 $T=1793880 2448880 1 0 $X=1793878 $Y=2443440
X44 5223 2 5132 4 5281 NAND2X1 $T=1803120 2509360 1 0 $X=1803118 $Y=2503920
X45 5261 2 5235 4 5236 NAND2X1 $T=1810380 2489200 1 180 $X=1808400 $Y=2488798
X46 5257 2 5251 4 5283 NAND2X1 $T=1817640 2509360 0 0 $X=1817638 $Y=2508958
X47 5321 2 5331 4 5303 NAND2X1 $T=1830180 2509360 0 0 $X=1830178 $Y=2508958
X48 5335 2 5333 4 5313 NAND2X1 $T=1832160 2529520 1 180 $X=1830180 $Y=2529118
X49 5333 2 5376 4 5377 NAND2X1 $T=1846020 2529520 1 0 $X=1846018 $Y=2524080
X50 5364 2 5408 4 5332 NAND2X1 $T=1848660 2499280 0 0 $X=1848658 $Y=2498878
X51 174 2 169 4 5407 NAND2X1 $T=1851300 2438800 1 0 $X=1851298 $Y=2433360
X52 141 2 5449 4 5444 NAND2X1 $T=1861860 2489200 0 0 $X=1861858 $Y=2488798
X53 141 2 5453 4 5448 NAND2X1 $T=1867140 2489200 0 0 $X=1867138 $Y=2488798
X54 5505 2 4703 4 5514 NAND2X1 $T=1879020 2458960 1 180 $X=1877040 $Y=2458558
X55 5281 2 5512 4 5511 NAND2X1 $T=1877700 2519440 0 0 $X=1877698 $Y=2519038
X56 5300 2 5331 4 5552 NAND2X1 $T=1885620 2499280 1 0 $X=1885618 $Y=2493840
X57 5331 2 5549 4 5559 NAND2X1 $T=1890240 2519440 1 0 $X=1890238 $Y=2514000
X58 5581 2 4937 4 5571 NAND2X1 $T=1894860 2469040 0 180 $X=1892880 $Y=2463600
X59 5533 2 5314 4 5621 NAND2X1 $T=1900800 2448880 1 0 $X=1900798 $Y=2443440
X60 5634 2 4907 4 5650 NAND2X1 $T=1908720 2479120 1 0 $X=1908718 $Y=2473680
X61 5686 2 196 4 5733 NAND2X1 $T=1927200 2489200 0 0 $X=1927198 $Y=2488798
X62 5768 2 5732 4 5800 NAND2X1 $T=1946340 2428720 1 0 $X=1946338 $Y=2423280
X63 5733 2 5802 4 5808 NAND2X1 $T=1950960 2479120 0 0 $X=1950958 $Y=2478718
X64 5830 2 5714 4 5752 NAND2X1 $T=1960200 2448880 1 0 $X=1960198 $Y=2443440
X65 5487 2 5106 4 5841 NAND2X1 $T=1966140 2469040 0 180 $X=1964160 $Y=2463600
X66 5443 2 202 4 5899 NAND2X1 $T=1981980 2428720 1 0 $X=1981978 $Y=2423280
X67 222 2 219 4 6569 NAND2X1 $T=2179980 2418640 0 180 $X=2178000 $Y=2413200
X68 6569 2 220 4 6555 NAND2X1 $T=2180640 2418640 0 0 $X=2180638 $Y=2418238
X69 2768 4 2 46 2840 NOR2X4 $T=1147080 2418640 0 180 $X=1142460 $Y=2413200
X70 3690 4 2 3696 3632 NOR2X4 $T=1390620 2489200 1 180 $X=1386000 $Y=2488798
X71 4190 4 2 4185 4071 NOR2X4 $T=1508760 2539600 1 0 $X=1508758 $Y=2534160
X72 3589 2 3605 3612 4 NAND2BX1 $T=1366200 2469040 1 180 $X=1363560 $Y=2468638
X73 3632 2 3631 3574 4 NAND2BX1 $T=1369500 2489200 1 180 $X=1366860 $Y=2488798
X74 94 2 91 3921 4 NAND2BX1 $T=1450020 2458960 1 180 $X=1447380 $Y=2458558
X75 3972 2 3971 3930 4 NAND2BX1 $T=1453320 2549680 0 180 $X=1450680 $Y=2544240
X76 3973 2 3934 3990 4 NAND2BX1 $T=1453320 2479120 1 0 $X=1453318 $Y=2473680
X77 4071 2 4051 4050 4 NAND2BX1 $T=1474440 2539600 1 180 $X=1471800 $Y=2539198
X78 4189 2 4192 4174 4 NAND2BX1 $T=1512060 2428720 0 180 $X=1509420 $Y=2423280
X79 4358 2 4296 4282 4 NAND2BX1 $T=1547700 2479120 0 180 $X=1545060 $Y=2473680
X80 4727 2 4725 4421 4 NAND2BX1 $T=1659900 2569840 0 180 $X=1657260 $Y=2564400
X81 4776 2 4795 165 4 NAND2BX1 $T=1681020 2569840 0 180 $X=1678380 $Y=2564400
X82 170 2 173 4938 4 NAND2BX1 $T=1717320 2428720 0 0 $X=1717318 $Y=2428318
X83 5154 2 5233 5177 4 NAND2BX1 $T=1806420 2438800 1 180 $X=1803780 $Y=2438398
X84 5103 2 5128 5274 4 NAND2BX1 $T=1813020 2438800 1 0 $X=1813018 $Y=2433360
X85 5381 2 5364 5297 4 NAND2BX1 $T=1843380 2499280 1 180 $X=1840740 $Y=2498878
X86 5410 2 5381 5450 4 NAND2BX1 $T=1853940 2499280 0 0 $X=1853938 $Y=2498878
X87 5622 2 5571 5623 4 NAND2BX1 $T=1900800 2458960 0 0 $X=1900798 $Y=2458558
X88 217 2 216 6479 4 NAND2BX1 $T=2162820 2418640 1 180 $X=2160180 $Y=2418238
X89 3588 3585 2 3575 4 3583 OAI21X1 $T=1356960 2529520 0 180 $X=1353660 $Y=2524080
X90 3590 3585 2 3587 4 3586 OAI21X1 $T=1358280 2509360 0 180 $X=1354980 $Y=2503920
X91 3624 3713 2 3772 4 3715 OAI21X1 $T=1401180 2519440 1 0 $X=1401178 $Y=2514000
X92 3902 3585 2 3839 4 3900 OAI21X1 $T=1440780 2539600 0 180 $X=1437480 $Y=2534160
X93 4106 4081 2 4109 4 4145 OAI21X1 $T=1488300 2489200 0 0 $X=1488298 $Y=2488798
X94 4406 4269 2 4396 4 4364 OAI21X1 $T=1570140 2529520 1 180 $X=1566840 $Y=2529118
X95 136 4269 2 4468 4 134 OAI21X1 $T=1591260 2569840 1 180 $X=1587960 $Y=2569438
X96 4547 4468 2 4604 4 4579 OAI21X1 $T=1624260 2559760 0 0 $X=1624258 $Y=2559358
X97 4727 161 2 4725 4 4661 OAI21X1 $T=1657260 2569840 0 0 $X=1657258 $Y=2569438
X98 5090 4595 2 5088 4 5129 OAI21X1 $T=1779360 2529520 0 180 $X=1776060 $Y=2524080
X99 5103 4290 2 5128 4 5176 OAI21X1 $T=1797180 2438800 1 0 $X=1797178 $Y=2433360
X100 5514 5622 2 5571 4 5574 OAI21X1 $T=1898160 2458960 1 180 $X=1894860 $Y=2458558
X101 5621 4290 2 5585 4 5584 OAI21X1 $T=1901460 2438800 1 180 $X=1898160 $Y=2438398
X102 217 6460 2 216 4 6554 OAI21X1 $T=2165460 2428720 1 0 $X=2165458 $Y=2423280
X103 216 221 2 6569 4 6583 OAI21X1 $T=2182620 2418640 0 0 $X=2182618 $Y=2418238
X104 67 2 54 68 4 3405 OAI21XL $T=1293600 2418640 1 0 $X=1293598 $Y=2413200
X105 3540 2 3604 3593 4 3645 OAI21XL $T=1359600 2428720 0 0 $X=1359598 $Y=2428318
X106 3789 2 3769 3770 4 3806 OAI21XL $T=1409100 2469040 1 0 $X=1409098 $Y=2463600
X107 3660 2 3585 3716 4 3865 OAI21XL $T=1424940 2519440 1 0 $X=1424938 $Y=2514000
X108 3770 2 3858 3874 4 3857 OAI21XL $T=1428900 2458960 0 180 $X=1426260 $Y=2453520
X109 3973 2 3864 3934 4 3922 OAI21XL $T=1449360 2479120 0 180 $X=1446720 $Y=2473680
X110 4109 2 4111 4170 4 4070 OAI21XL $T=1491600 2469040 0 180 $X=1488960 $Y=2463600
X111 4192 2 4249 4220 4 4240 OAI21XL $T=1526580 2428720 0 0 $X=1526578 $Y=2428318
X112 4296 2 4363 4403 4 4404 OAI21XL $T=1567500 2499280 1 0 $X=1567498 $Y=2493840
X113 4446 2 4423 4475 4 4474 OAI21XL $T=1593240 2529520 1 180 $X=1590600 $Y=2529118
X114 4678 2 4776 4795 4 4710 OAI21XL $T=1679700 2559760 1 180 $X=1677060 $Y=2559358
X115 170 2 116 4743 4 4920 OAI21XL $T=1710720 2438800 1 0 $X=1710718 $Y=2433360
X116 4938 2 116 4939 4 4971 OAI21XL $T=1718640 2438800 0 0 $X=1718638 $Y=2438398
X117 5088 2 5117 5116 4 5115 OAI21XL $T=1774740 2519440 0 180 $X=1772100 $Y=2514000
X118 5255 2 4595 5236 4 180 OAI21XL $T=1810380 2479120 1 180 $X=1807740 $Y=2478718
X119 5259 2 4595 5250 4 181 OAI21XL $T=1811700 2458960 1 180 $X=1809060 $Y=2458558
X120 5313 2 5258 5306 4 5235 OAI21XL $T=1826220 2529520 0 180 $X=1823580 $Y=2524080
X121 5332 2 5300 5297 4 5336 OAI21XL $T=1839420 2509360 0 180 $X=1836780 $Y=2503920
X122 5350 2 4595 5349 4 184 OAI21XL $T=1840740 2438800 0 180 $X=1838100 $Y=2433360
X123 5283 2 4595 5263 4 187 OAI21XL $T=1842060 2448880 1 0 $X=1842058 $Y=2443440
X124 5410 2 5300 5381 4 5412 OAI21XL $T=1851300 2509360 0 0 $X=1851298 $Y=2508958
X125 5317 2 4595 5414 4 5422 OAI21XL $T=1852620 2458960 0 0 $X=1852618 $Y=2458558
X126 5413 2 4595 5409 4 188 OAI21XL $T=1853940 2448880 1 0 $X=1853938 $Y=2443440
X127 5444 2 4595 5448 4 5457 OAI21XL $T=1861200 2489200 1 0 $X=1861198 $Y=2483760
X128 5258 2 5377 5445 4 5453 OAI21XL $T=1861200 2519440 0 0 $X=1861198 $Y=2519038
X129 5485 2 4595 5455 4 5488 OAI21XL $T=1870440 2499280 0 0 $X=1870438 $Y=2498878
X130 5277 2 4595 5258 4 5526 OAI21XL $T=1882320 2519440 0 0 $X=1882318 $Y=2519038
X131 5559 2 4595 5541 4 5561 OAI21XL $T=1891560 2509360 0 0 $X=1891558 $Y=2508958
X132 5806 2 193 5805 4 5801 OAI21XL $T=1953600 2448880 0 180 $X=1950960 $Y=2443440
X133 5841 2 5900 5899 4 5858 OAI21XL $T=1987920 2458960 1 0 $X=1987918 $Y=2453520
X134 142 116 4318 2 4 XOR2X4 $T=1613700 2418640 0 180 $X=1602480 $Y=2413200
X135 174 224 225 2 4 XOR2X4 $T=2282280 2428720 0 0 $X=2282278 $Y=2428318
X136 46 2 4 47 INVX1 $T=1151040 2418640 1 0 $X=1151038 $Y=2413200
X137 3623 2 4 3590 INVX1 $T=1364220 2509360 0 180 $X=1362900 $Y=2503920
X138 3646 2 4 3587 INVX1 $T=1371480 2509360 0 180 $X=1370160 $Y=2503920
X139 3624 2 4 3614 INVX1 $T=1374120 2529520 0 180 $X=1372800 $Y=2524080
X140 3663 2 4 3613 INVX1 $T=1379400 2529520 1 0 $X=1379398 $Y=2524080
X141 83 2 4 3769 INVX1 $T=1410420 2479120 0 0 $X=1410418 $Y=2478718
X142 3876 2 4 3841 INVX1 $T=1424280 2539600 1 180 $X=1422960 $Y=2539198
X143 3875 2 4 3878 INVX1 $T=1430880 2539600 1 0 $X=1430878 $Y=2534160
X144 3716 2 4 4028 INVX1 $T=1472460 2539600 1 0 $X=1472458 $Y=2534160
X145 3899 2 4 4123 INVX1 $T=1490280 2519440 0 0 $X=1490278 $Y=2519038
X146 4377 2 4 4308 INVX1 $T=1557600 2519440 1 180 $X=1556280 $Y=2519038
X147 4295 2 4 4429 INVX1 $T=1576740 2519440 1 0 $X=1576738 $Y=2514000
X148 4446 2 4 4405 INVX1 $T=1581360 2519440 0 180 $X=1580040 $Y=2514000
X149 4269 2 4 144 INVX1 $T=1589940 2569840 1 0 $X=1589938 $Y=2564400
X150 4531 2 4 4407 INVX1 $T=1607100 2529520 0 180 $X=1605780 $Y=2524080
X151 4468 2 4 148 INVX1 $T=1626900 2569840 0 0 $X=1626898 $Y=2569438
X152 4646 2 4 4556 INVX1 $T=1633500 2559760 1 180 $X=1632180 $Y=2559358
X153 4640 2 4 4658 INVX1 $T=1638120 2549680 0 0 $X=1638118 $Y=2549278
X154 167 2 4 4757 INVX1 $T=1680360 2418640 0 180 $X=1679040 $Y=2413200
X155 4743 2 4 4972 INVX1 $T=1729200 2438800 0 0 $X=1729198 $Y=2438398
X156 5177 2 4 5173 INVX1 $T=1797840 2438800 1 180 $X=1796520 $Y=2438398
X157 5115 2 4 5258 INVX1 $T=1798500 2529520 1 0 $X=1798498 $Y=2524080
X158 5251 2 4 5277 INVX1 $T=1809720 2519440 0 0 $X=1809718 $Y=2519038
X159 5321 2 4 5302 INVX1 $T=1826880 2509360 0 180 $X=1825560 $Y=2503920
X160 5280 2 4 5317 INVX1 $T=1826880 2458960 0 0 $X=1826878 $Y=2458558
X161 5283 2 4 5353 INVX1 $T=1833480 2448880 0 0 $X=1833478 $Y=2448478
X162 5263 2 4 5318 INVX1 $T=1834800 2448880 0 180 $X=1833480 $Y=2443440
X163 146 2 4 183 INVX1 $T=1836120 2418640 1 0 $X=1836118 $Y=2413200
X164 5235 2 4 5414 INVX1 $T=1836120 2469040 1 0 $X=1836118 $Y=2463600
X165 5281 2 4 5411 INVX1 $T=1838760 2519440 0 0 $X=1838758 $Y=2519038
X166 5253 2 4 5333 INVX1 $T=1838760 2529520 0 0 $X=1838758 $Y=2529118
X167 5331 2 4 5347 INVX1 $T=1846680 2519440 1 0 $X=1846678 $Y=2514000
X168 5410 2 4 5408 INVX1 $T=1850640 2499280 0 180 $X=1849320 $Y=2493840
X169 5453 2 4 5455 INVX1 $T=1863180 2499280 0 0 $X=1863178 $Y=2498878
X170 5449 2 4 5485 INVX1 $T=1863180 2509360 1 0 $X=1863178 $Y=2503920
X171 5300 2 4 5540 INVX1 $T=1877700 2509360 1 0 $X=1877698 $Y=2503920
X172 5260 2 4 5513 INVX1 $T=1881660 2438800 1 180 $X=1880340 $Y=2438398
X173 5314 2 4 5507 INVX1 $T=1881660 2448880 0 180 $X=1880340 $Y=2443440
X174 5529 2 4 5533 INVX1 $T=1885620 2458960 1 0 $X=1885618 $Y=2453520
X175 4595 2 4 5567 INVX1 $T=1898820 2519440 0 0 $X=1898818 $Y=2519038
X176 5666 2 4 5701 INVX1 $T=1929840 2469040 1 0 $X=1929838 $Y=2463600
X177 5752 2 4 5768 INVX1 $T=1941720 2428720 0 180 $X=1940400 $Y=2423280
X178 5653 2 4 5803 INVX1 $T=1945680 2438800 1 0 $X=1945678 $Y=2433360
X179 213 2 4 6395 INVX1 $T=2121240 2418640 0 0 $X=2121238 $Y=2418238
X180 42 41 4 43 2702 2 AOI21X2 $T=1097580 2418640 1 0 $X=1097578 $Y=2413200
X181 52 2840 4 2781 50 2 AOI21X2 $T=1186680 2418640 1 180 $X=1182060 $Y=2418238
X182 3122 2781 4 3141 3143 2 AOI21X2 $T=1221000 2418640 0 0 $X=1220998 $Y=2418238
X183 3438 52 4 3405 69 2 AOI21X2 $T=1304160 2418640 0 180 $X=1299540 $Y=2413200
X184 79 78 4 77 3504 2 AOI21X2 $T=1360920 2418640 0 180 $X=1356300 $Y=2413200
X185 3840 83 4 3857 3864 2 AOI21X2 $T=1425600 2479120 1 0 $X=1425598 $Y=2473680
X186 4065 3986 4 4070 4035 2 AOI21X2 $T=1477080 2469040 0 0 $X=1477078 $Y=2468638
X187 4117 3996 4 4130 4139 2 AOI21X2 $T=1492260 2549680 0 0 $X=1492258 $Y=2549278
X188 4473 4429 4 4474 4468 2 AOI21X2 $T=1587300 2539600 0 0 $X=1587298 $Y=2539198
X189 4 61 59 3122 2 NOR2X1 $T=1250700 2418640 0 180 $X=1248720 $Y=2413200
X190 4 59 56 64 2 NOR2X1 $T=1259940 2418640 1 0 $X=1259938 $Y=2413200
X191 4 65 56 66 2 NOR2X1 $T=1287660 2418640 1 0 $X=1287658 $Y=2413200
X192 4 67 56 3438 2 NOR2X1 $T=1307460 2418640 1 0 $X=1307458 $Y=2413200
X193 4 3530 3604 3630 2 NOR2X1 $T=1362240 2438800 1 0 $X=1362238 $Y=2433360
X194 4 3614 3608 3575 2 NOR2X1 $T=1364220 2529520 0 180 $X=1362240 $Y=2524080
X195 4 3626 80 3589 2 NOR2X1 $T=1366860 2489200 0 180 $X=1364880 $Y=2483760
X196 4 3632 3589 3623 2 NOR2X1 $T=1367520 2499280 1 180 $X=1365540 $Y=2498878
X197 4 3680 81 3530 2 NOR2X1 $T=1375440 2428720 1 180 $X=1373460 $Y=2428318
X198 4 3803 3773 3663 2 NOR2X1 $T=1405800 2529520 0 180 $X=1403820 $Y=2524080
X199 4 85 84 3789 2 NOR2X1 $T=1421640 2438800 0 180 $X=1419660 $Y=2433360
X200 4 3789 3858 3840 2 NOR2X1 $T=1426920 2469040 1 0 $X=1426918 $Y=2463600
X201 4 90 3904 3875 2 NOR2X1 $T=1445400 2539600 0 0 $X=1445398 $Y=2539198
X202 4 95 93 3973 2 NOR2X1 $T=1455300 2438800 1 0 $X=1455298 $Y=2433360
X203 4 94 3973 4015 2 NOR2X1 $T=1457940 2458960 0 0 $X=1457938 $Y=2458558
X204 4 4111 4106 4065 2 NOR2X1 $T=1490280 2479120 0 180 $X=1488300 $Y=2473680
X205 4 103 102 4106 2 NOR2X1 $T=1490940 2458960 0 180 $X=1488960 $Y=2453520
X206 4 4120 4123 4146 2 NOR2X1 $T=1492920 2519440 1 0 $X=1492918 $Y=2514000
X207 4 106 107 4111 2 NOR2X1 $T=1502160 2469040 1 0 $X=1502158 $Y=2463600
X208 4 4249 4189 111 2 NOR2X1 $T=1539120 2428720 0 0 $X=1539118 $Y=2428318
X209 4 4343 4319 4249 2 NOR2X1 $T=1551660 2428720 1 180 $X=1549680 $Y=2428318
X210 4 4395 4361 4358 2 NOR2X1 $T=1559580 2479120 0 180 $X=1557600 $Y=2473680
X211 4 4358 4363 4377 2 NOR2X1 $T=1560900 2489200 0 0 $X=1560898 $Y=2488798
X212 4 4412 4420 4363 2 NOR2X1 $T=1576080 2489200 1 180 $X=1574100 $Y=2488798
X213 4 4497 4488 4531 2 NOR2X1 $T=1600500 2519440 1 0 $X=1600498 $Y=2514000
X214 4 4423 4531 4473 2 NOR2X1 $T=1602480 2529520 0 0 $X=1602478 $Y=2529118
X215 4 4547 136 4560 2 NOR2X1 $T=1607760 2559760 0 0 $X=1607758 $Y=2559358
X216 4 4640 4556 149 2 NOR2X1 $T=1633500 2569840 1 180 $X=1631520 $Y=2569438
X217 4 4739 4704 4727 2 NOR2X1 $T=1653960 2549680 1 180 $X=1651980 $Y=2549278
X218 4 4776 4640 4708 2 NOR2X1 $T=1666500 2559760 1 180 $X=1664520 $Y=2559358
X219 4 4890 4840 4776 2 NOR2X1 $T=1700820 2549680 1 180 $X=1698840 $Y=2549278
X220 4 5072 4954 5090 2 NOR2X1 $T=1758240 2529520 1 0 $X=1758238 $Y=2524080
X221 4 5102 177 5103 2 NOR2X1 $T=1764840 2438800 1 0 $X=1764838 $Y=2433360
X222 4 5085 5105 5117 2 NOR2X1 $T=1780680 2509360 0 0 $X=1780678 $Y=2508958
X223 4 5157 178 5154 2 NOR2X1 $T=1789920 2438800 1 180 $X=1787940 $Y=2438398
X224 4 5117 5090 5251 2 NOR2X1 $T=1799160 2519440 0 0 $X=1799158 $Y=2519038
X225 4 5223 5132 5253 2 NOR2X1 $T=1803120 2509360 0 0 $X=1803118 $Y=2508958
X226 4 5253 5303 5257 2 NOR2X1 $T=1824240 2509360 1 180 $X=1822260 $Y=2508958
X227 4 5313 5277 5280 2 NOR2X1 $T=1828860 2519440 0 180 $X=1826880 $Y=2514000
X228 4 5296 5332 5321 2 NOR2X1 $T=1830180 2499280 0 0 $X=1830178 $Y=2498878
X229 4 5332 5347 5335 2 NOR2X1 $T=1837440 2519440 0 180 $X=1835460 $Y=2514000
X230 4 183 186 5364 2 NOR2X1 $T=1840740 2479120 1 0 $X=1840738 $Y=2473680
X231 4 132 5366 5410 2 NOR2X1 $T=1851300 2489200 1 0 $X=1851298 $Y=2483760
X232 4 5410 5347 5376 2 NOR2X1 $T=1853280 2519440 0 180 $X=1851300 $Y=2514000
X233 4 5377 5277 5449 2 NOR2X1 $T=1859220 2519440 1 0 $X=1859218 $Y=2514000
X234 4 5253 5277 5549 2 NOR2X1 $T=1875060 2519440 1 0 $X=1875058 $Y=2514000
X235 4 5505 4703 5529 2 NOR2X1 $T=1882320 2458960 0 0 $X=1882318 $Y=2458558
X236 4 5634 4907 5666 2 NOR2X1 $T=1913340 2479120 1 0 $X=1913338 $Y=2473680
X237 4 5487 5106 5831 2 NOR2X1 $T=1962840 2458960 1 180 $X=1960860 $Y=2458558
X238 4 5443 202 5900 2 NOR2X1 $T=1983960 2428720 1 0 $X=1983958 $Y=2423280
X239 4 217 221 6570 2 NOR2X1 $T=2180640 2438800 1 0 $X=2180638 $Y=2433360
X240 4 222 219 221 2 NOR2X1 $T=2187900 2418640 1 0 $X=2187898 $Y=2413200
X241 3712 82 2 4 3604 NOR2X2 $T=1391280 2438800 0 180 $X=1387980 $Y=2433360
X242 3713 3663 2 4 3698 NOR2X2 $T=1391940 2529520 1 0 $X=1391938 $Y=2524080
X243 87 86 2 4 3858 NOR2X2 $T=1429560 2418640 0 0 $X=1429558 $Y=2418238
X244 3974 3995 2 4 3713 NOR2X2 $T=1455300 2519440 0 180 $X=1452000 $Y=2514000
X245 3972 3875 2 4 4012 NOR2X2 $T=1457280 2539600 0 0 $X=1457278 $Y=2539198
X246 4043 4033 2 4 3972 NOR2X2 $T=1469160 2549680 1 0 $X=1469158 $Y=2544240
X247 4071 4188 2 4 4117 NOR2X2 $T=1511400 2559760 0 180 $X=1508100 $Y=2554320
X248 4318 120 2 4 4188 NOR2X2 $T=1545720 2549680 1 180 $X=1542420 $Y=2549278
X249 4312 119 2 4 4189 NOR2X2 $T=1547700 2418640 1 0 $X=1547698 $Y=2413200
X250 4568 4559 2 4 4423 NOR2X2 $T=1615020 2529520 0 0 $X=1615018 $Y=2529118
X251 139 4727 2 4 4646 NOR2X2 $T=1655280 2569840 1 180 $X=1651980 $Y=2569438
X252 4792 4774 2 4 4640 NOR2X2 $T=1675080 2549680 0 180 $X=1671780 $Y=2544240
X253 5103 5154 2 4 5314 NOR2X2 $T=1818300 2438800 0 0 $X=1818298 $Y=2438398
X254 4937 5581 2 4 5622 NOR2X2 $T=1902780 2469040 0 0 $X=1902778 $Y=2468638
X255 5529 5622 2 4 5632 NOR2X2 $T=1905420 2458960 0 0 $X=1905418 $Y=2458558
X256 196 5686 2 4 5697 NOR2X2 $T=1929180 2489200 0 180 $X=1925880 $Y=2483760
X257 5666 5697 2 4 5714 NOR2X2 $T=1933140 2479120 0 180 $X=1929840 $Y=2473680
X258 5653 5752 2 4 197 NOR2X2 $T=1941060 2428720 1 180 $X=1937760 $Y=2428318
X259 5831 5900 2 4 5830 NOR2X2 $T=1983300 2458960 0 180 $X=1980000 $Y=2453520
X260 167 152 2 4 4810 OR2XL $T=1687620 2418640 0 180 $X=1684980 $Y=2413200
X261 3913 3971 3996 2 4 NAND2X2 $T=1462560 2549680 1 180 $X=1459260 $Y=2549278
X262 4577 4602 4582 2 4 NAND2X2 $T=1620960 2569840 1 180 $X=1617660 $Y=2569438
X263 5314 5632 5653 2 4 NAND2X2 $T=1908720 2448880 1 0 $X=1908718 $Y=2443440
X264 5800 5777 199 2 4 NAND2X2 $T=1951620 2418640 0 180 $X=1948320 $Y=2413200
X265 3698 4 3646 3715 2 3716 AOI21X4 $T=1389960 2519440 1 0 $X=1389958 $Y=2514000
X266 4560 4 144 4579 2 4595 AOI21X4 $T=1613700 2559760 0 0 $X=1613698 $Y=2559358
X267 5632 4 5260 5574 2 5637 AOI21X4 $T=1904100 2458960 1 0 $X=1904098 $Y=2453520
X268 6570 4 6504 6583 2 223 AOI21X4 $T=2180640 2428720 1 0 $X=2180638 $Y=2423280
X269 3613 4 3646 2 3608 AND2X2 $T=1364220 2509360 1 180 $X=1361580 $Y=2508958
X270 3630 4 78 2 3654 AND2X2 $T=1368180 2418640 1 0 $X=1368178 $Y=2413200
X271 4012 4 3899 2 4018 AND2X2 $T=1461240 2529520 0 0 $X=1461238 $Y=2529118
X272 4079 4 3899 2 4093 AND2X2 $T=1482360 2529520 1 0 $X=1482358 $Y=2524080
X273 162 4 156 2 5261 AND2X2 $T=1806420 2479120 1 0 $X=1806418 $Y=2473680
X274 5701 4 5650 2 5682 AND2X2 $T=1925880 2469040 0 180 $X=1923240 $Y=2463600
X275 5824 4 5803 2 5804 AND2X2 $T=1955580 2438800 0 180 $X=1952940 $Y=2433360
X276 211 4 209 2 6377 AND2X2 $T=2113320 2428720 1 0 $X=2113318 $Y=2423280
X277 42 2 44 4 2768 NAND2X4 $T=1108800 2418640 1 0 $X=1108798 $Y=2413200
X278 3972 3876 2 4 3913 OR2X2 $T=1446060 2549680 1 180 $X=1443420 $Y=2549278
X279 5158 5315 2 4 5331 OR2X2 $T=1827540 2489200 0 0 $X=1827538 $Y=2488798
X280 5263 5407 2 4 5409 OR2X2 $T=1848660 2448880 1 0 $X=1848658 $Y=2443440
X281 5283 5407 2 4 5413 OR2X2 $T=1851300 2458960 1 0 $X=1851298 $Y=2453520
X282 5258 5253 2 4 5512 OR2X2 $T=1871760 2519440 0 0 $X=1871758 $Y=2519038
X283 5653 5666 2 4 5723 OR2X2 $T=1924560 2448880 0 0 $X=1924558 $Y=2448478
X284 5697 5650 2 4 5802 OR2X2 $T=1950300 2479120 1 0 $X=1950298 $Y=2473680
X285 4678 2 4 4658 4593 NAND2XL $T=1644060 2549680 0 180 $X=1642080 $Y=2544240
X286 4757 2 4 160 4773 NAND2XL $T=1673760 2418640 1 0 $X=1673758 $Y=2413200
X287 5085 2 4 5105 5116 NAND2XL $T=1770120 2509360 0 0 $X=1770118 $Y=2508958
X288 156 2 4 5235 5250 NAND2XL $T=1806420 2469040 1 0 $X=1806418 $Y=2463600
X289 166 2 4 5261 5296 NAND2XL $T=1815000 2499280 1 0 $X=1814998 $Y=2493840
X290 156 2 4 5280 5259 NAND2XL $T=1816980 2458960 1 180 $X=1815000 $Y=2458558
X291 5261 2 4 5280 5255 NAND2XL $T=1817640 2479120 0 0 $X=1817638 $Y=2478718
X292 5315 2 4 5158 5300 NAND2XL $T=1824240 2489200 1 180 $X=1822260 $Y=2488798
X293 169 2 4 5318 5349 NAND2XL $T=1827540 2438800 0 0 $X=1827538 $Y=2438398
X294 169 2 4 5353 5350 NAND2XL $T=1841400 2458960 0 180 $X=1839420 $Y=2453520
X295 132 2 4 5366 5381 NAND2XL $T=1846020 2489200 1 0 $X=1846018 $Y=2483760
X296 5514 2 4 5533 5490 NAND2XL $T=1881000 2458960 0 180 $X=1879020 $Y=2453520
X297 5714 2 4 5803 5806 NAND2XL $T=1958220 2448880 0 180 $X=1956240 $Y=2443440
X298 213 2 4 211 214 NAND2XL $T=2125860 2418640 0 0 $X=2125858 $Y=2418238
X299 4266 4269 2 4 INVX4 $T=1537800 2469040 0 180 $X=1535160 $Y=2463600
X300 3630 77 4 3645 3662 2 AOI21X1 $T=1369500 2428720 1 0 $X=1369498 $Y=2423280
X301 4012 4028 4 3996 4046 2 AOI21X1 $T=1465200 2539600 1 0 $X=1465198 $Y=2534160
X302 4028 4079 4 4080 4105 2 AOI21X1 $T=1479720 2539600 1 0 $X=1479718 $Y=2534160
X303 3676 4146 4 4172 4202 2 AOI21X1 $T=1500840 2519440 1 0 $X=1500838 $Y=2514000
X304 112 111 4 4240 4239 2 AOI21X1 $T=1527240 2418640 1 180 $X=1524600 $Y=2418238
X305 4407 4404 4 4405 4396 2 AOI21X1 $T=1571460 2519440 1 180 $X=1568820 $Y=2519038
X306 4646 148 4 4661 4602 2 AOI21X1 $T=1642080 2569840 0 0 $X=1642078 $Y=2569438
X307 4661 4708 4 4710 4604 2 AOI21X1 $T=1654620 2559760 0 0 $X=1654618 $Y=2559358
X308 173 4972 4 175 4939 2 AOI21X1 $T=1729200 2438800 1 0 $X=1729198 $Y=2433360
X309 5256 5257 4 5262 5263 2 AOI21X1 $T=1811700 2509360 0 0 $X=1811698 $Y=2508958
X310 5376 5411 4 5412 5445 2 AOI21X1 $T=1851300 2529520 1 0 $X=1851298 $Y=2524080
X311 5701 5732 4 5734 5731 2 AOI21X1 $T=1937760 2469040 1 0 $X=1937758 $Y=2463600
X312 5732 5824 4 5829 5807 2 AOI21X1 $T=1958880 2438800 1 0 $X=1958878 $Y=2433360
X313 5808 5830 4 5858 5777 2 AOI21X1 $T=1968780 2458960 1 0 $X=1968778 $Y=2453520
X314 212 211 4 6395 6378 2 AOI21X1 $T=2123220 2428720 1 0 $X=2123218 $Y=2423280
X315 3530 3504 2 3540 4 3503 OAI21X2 $T=1345740 2438800 1 0 $X=1345738 $Y=2433360
X316 3589 3585 2 3605 4 3573 OAI21X2 $T=1356300 2479120 1 0 $X=1356298 $Y=2473680
X317 3657 3632 2 3631 4 3646 OAI21X2 $T=1379400 2499280 0 180 $X=1374120 $Y=2493840
X318 3934 94 2 91 4 3986 OAI21X2 $T=1455960 2448880 1 180 $X=1450680 $Y=2448478
X319 4030 3864 2 4035 4 4048 OAI21X2 $T=1466520 2469040 0 0 $X=1466518 $Y=2468638
X320 4120 3716 2 4139 4 4172 OAI21X2 $T=1493580 2529520 1 0 $X=1493578 $Y=2524080
X321 4189 108 2 4192 4 4129 OAI21X2 $T=1508100 2428720 0 0 $X=1508098 $Y=2428318
X322 4051 4188 2 4203 4 4130 OAI21X2 $T=1508100 2549680 0 0 $X=1508098 $Y=2549278
X323 4308 4269 2 4295 4 4268 OAI21X2 $T=1549680 2519440 1 180 $X=1544400 $Y=2519038
X324 4358 4269 2 4296 4 4317 OAI21X2 $T=1550340 2489200 1 180 $X=1545060 $Y=2488798
X325 4269 129 2 4454 4 4424 OAI21X2 $T=1579380 2569840 0 0 $X=1579378 $Y=2569438
X326 5128 5154 2 5233 4 5260 OAI21X2 $T=1814340 2438800 1 180 $X=1809060 $Y=2438398
X327 5507 4290 2 5513 4 5486 OAI21X2 $T=1877040 2438800 1 0 $X=1877038 $Y=2433360
X328 5653 193 2 5637 4 5684 OAI21X2 $T=1916640 2438800 1 180 $X=1911360 $Y=2438398
X329 5723 193 2 5731 4 5721 OAI21X2 $T=1934460 2458960 1 0 $X=1934458 $Y=2453520
X330 3505 3503 71 2 4 XNOR2X4 $T=1338480 2438800 1 180 $X=1327260 $Y=2438398
X331 4593 4582 4190 2 4 XNOR2X4 $T=1623600 2549680 0 180 $X=1612380 $Y=2544240
X332 45 2 2768 2702 4 2781 OAI21X4 $T=1123980 2418640 0 180 $X=1116720 $Y=2413200
X333 3120 2 57 3143 4 58 OAI21X4 $T=1221000 2418640 1 0 $X=1220998 $Y=2413200
X334 3515 3504 4 2 72 XOR2X2 $T=1339140 2428720 1 180 $X=1332540 $Y=2428318
X335 3584 3583 4 2 74 XOR2X2 $T=1357620 2519440 0 180 $X=1351020 $Y=2514000
X336 3612 3585 4 2 75 XOR2X2 $T=1364220 2458960 1 180 $X=1357620 $Y=2458558
X337 4087 4081 4 2 4043 XOR2X2 $T=1484340 2499280 0 180 $X=1477740 $Y=2493840
X338 4174 108 4 2 3680 XOR2X2 $T=1504800 2428720 0 180 $X=1498200 $Y=2423280
X339 4282 4269 4 2 3626 XOR2X2 $T=1540440 2479120 0 180 $X=1533840 $Y=2473680
X340 4320 4317 4 2 3690 XOR2X2 $T=1552320 2499280 1 180 $X=1545720 $Y=2498878
X341 4365 4364 4 2 3995 XOR2X2 $T=1561560 2529520 1 180 $X=1554960 $Y=2529118
X342 5173 5176 4 2 179 XOR2X2 $T=1793880 2428720 1 0 $X=1793878 $Y=2423280
X343 5274 4290 4 2 182 XOR2X2 $T=1814340 2428720 1 0 $X=1814338 $Y=2423280
X344 156 190 4 2 192 XOR2X2 $T=1872420 2418640 1 0 $X=1872418 $Y=2413200
X345 5682 5684 4 2 195 XOR2X2 $T=1919940 2438800 1 0 $X=1919938 $Y=2433360
X346 6479 6460 4 2 215 XOR2X2 $T=2148300 2428720 0 180 $X=2141700 $Y=2423280
X347 2840 2 56 4 INVX2 $T=1210440 2418640 0 0 $X=1210438 $Y=2418238
X348 3660 2 3899 4 INVX2 $T=1437480 2519440 1 0 $X=1437478 $Y=2514000
X349 3864 2 3989 4 INVX2 $T=1461900 2479120 0 0 $X=1461898 $Y=2478718
X350 5637 2 5732 4 INVX2 $T=1956240 2458960 1 0 $X=1956238 $Y=2453520
X351 4071 4 2 4067 INVXL $T=1484340 2549680 1 180 $X=1483020 $Y=2549278
X352 5258 4 2 5256 INVXL $T=1812360 2529520 1 0 $X=1812358 $Y=2524080
X353 156 4 2 185 INVXL $T=1844040 2418640 1 0 $X=1844038 $Y=2413200
X354 5514 4 2 5564 INVXL $T=1890900 2458960 0 0 $X=1890898 $Y=2458558
X355 5511 4 2 5563 INVXL $T=1893540 2529520 0 0 $X=1893538 $Y=2529118
X356 5650 4 2 5734 INVXL $T=1941720 2469040 1 180 $X=1940400 $Y=2468638
X357 5714 4 2 5821 INVXL $T=1953600 2469040 1 0 $X=1953598 $Y=2463600
X358 5831 4 2 5871 INVXL $T=1982640 2458960 0 0 $X=1982638 $Y=2458558
X359 3574 3573 4 2 73 XNOR2X2 $T=1353000 2479120 0 180 $X=1345740 $Y=2473680
X360 4134 4129 4 2 3712 XNOR2X2 $T=1497540 2438800 0 180 $X=1490280 $Y=2433360
X361 4171 4145 4 2 4185 XNOR2X2 $T=1500180 2489200 0 0 $X=1500178 $Y=2488798
X362 4256 4223 4 2 115 XNOR2X2 $T=1528560 2539600 1 0 $X=1528558 $Y=2534160
X363 4270 4268 4 2 3803 XNOR2X2 $T=1537800 2529520 0 180 $X=1530540 $Y=2524080
X364 4421 4424 4 2 4033 XNOR2X2 $T=1578060 2569840 0 180 $X=1570800 $Y=2564400
X365 5144 5129 4 2 5157 XNOR2X2 $T=1783980 2529520 1 0 $X=1783978 $Y=2524080
X366 5552 5560 4 2 5581 XNOR2X2 $T=1890900 2499280 1 0 $X=1890898 $Y=2493840
X367 5623 5584 4 2 191 XNOR2X2 $T=1905420 2428720 1 180 $X=1898160 $Y=2428318
X368 5718 5721 4 2 198 XNOR2X2 $T=1931820 2448880 1 0 $X=1931818 $Y=2443440
X369 5870 5801 4 2 201 XNOR2X2 $T=1974060 2448880 1 0 $X=1974058 $Y=2443440
X370 6555 6554 4 2 218 XNOR2X2 $T=2175360 2418640 1 180 $X=2168100 $Y=2418238
X371 3768 3769 2 4 3696 XOR2X1 $T=1401180 2479120 0 180 $X=1395900 $Y=2473680
X372 3823 3806 2 4 3773 XOR2X1 $T=1417020 2469040 1 180 $X=1411740 $Y=2468638
X373 176 4971 2 4 5106 XOR2X1 $T=1739100 2438800 0 0 $X=1739098 $Y=2438398
X374 5086 4595 2 4 5102 XOR2X1 $T=1761540 2458960 0 0 $X=1761538 $Y=2458558
X375 3772 4 3713 3584 2 NOR2BX1 $T=1413060 2519440 0 180 $X=1410420 $Y=2514000
X376 3874 4 3858 3823 2 NOR2BX1 $T=1431540 2448880 0 180 $X=1428900 $Y=2443440
X377 4012 4 4071 4079 2 NOR2BX1 $T=1479720 2539600 0 0 $X=1479718 $Y=2539198
X378 4403 4 4363 4320 2 NOR2BX1 $T=1560900 2499280 0 180 $X=1558260 $Y=2493840
X379 4475 4 4423 4365 2 NOR2BX1 $T=1578720 2529520 1 180 $X=1576080 $Y=2529118
X380 5714 4 5831 5824 2 NOR2BX1 $T=1966140 2448880 1 0 $X=1966138 $Y=2443440
X381 131 127 123 4401 4 2 4383 ADDFX2 $T=1580700 2438800 0 180 $X=1566840 $Y=2433360
X382 4441 4440 4419 4412 4 2 4361 ADDFX2 $T=1584000 2469040 1 180 $X=1570140 $Y=2468638
X383 4535 4500 4501 4497 4 2 4420 ADDFX2 $T=1606440 2479120 1 180 $X=1592580 $Y=2478718
X384 130 141 128 4500 4 2 4419 ADDFX2 $T=1609080 2469040 1 180 $X=1595220 $Y=2468638
X385 137 123 128 4545 4 2 4535 ADDFX2 $T=1595880 2448880 1 0 $X=1595878 $Y=2443440
X386 4580 4581 4565 4559 4 2 4488 ADDFX2 $T=1624260 2499280 1 180 $X=1610400 $Y=2498878
X387 132 146 4591 4580 4 2 4501 ADDFX2 $T=1630860 2479120 0 180 $X=1617000 $Y=2473680
X388 143 130 132 4615 4 2 4581 ADDFX2 $T=1618980 2489200 1 0 $X=1618978 $Y=2483760
X389 4669 4706 4679 154 4 2 4568 ADDFX2 $T=1658580 2529520 0 180 $X=1644720 $Y=2524080
X390 147 128 141 4723 4 2 4706 ADDFX2 $T=1645380 2469040 0 0 $X=1645378 $Y=2468638
X391 141 156 4545 4669 4 2 4565 ADDFX2 $T=1659240 2499280 0 180 $X=1645380 $Y=2493840
X392 146 162 4615 4701 4 2 4679 ADDFX2 $T=1663200 2489200 0 180 $X=1649340 $Y=2483760
X393 4701 4707 4726 4739 4 2 163 ADDFX2 $T=1650660 2509360 0 0 $X=1650658 $Y=2508958
X394 158 132 146 4756 4 2 4707 ADDFX2 $T=1655940 2469040 1 0 $X=1655938 $Y=2463600
X395 156 166 4723 4772 4 2 4726 ADDFX2 $T=1684980 2499280 1 180 $X=1671120 $Y=2498878
X396 4772 4809 4789 4774 4 2 4704 ADDFX2 $T=1687620 2509360 0 180 $X=1673760 $Y=2503920
X397 162 169 4756 4836 4 2 4789 ADDFX2 $T=1704120 2479120 0 180 $X=1690260 $Y=2473680
X398 4836 4892 4844 4840 4 2 4792 ADDFX2 $T=1706100 2539600 0 180 $X=1692240 $Y=2534160
X399 172 141 156 4956 4 2 4809 ADDFX2 $T=1713360 2499280 1 0 $X=1713358 $Y=2493840
X400 166 174 4956 4952 4 2 4844 ADDFX2 $T=1733820 2509360 0 180 $X=1719960 $Y=2503920
X401 131 146 162 4982 4 2 4892 ADDFX2 $T=1720620 2479120 1 0 $X=1720618 $Y=2473680
X402 4989 4982 4952 4954 4 2 4890 ADDFX2 $T=1735140 2539600 0 180 $X=1721280 $Y=2534160
X403 166 169 5027 5022 4 2 4989 ADDFX2 $T=1755600 2499280 0 180 $X=1741740 $Y=2493840
X404 5022 5062 5073 5085 4 2 5072 ADDFX2 $T=1750320 2509360 1 0 $X=1750318 $Y=2503920
X405 169 174 5087 5075 4 2 5073 ADDFX2 $T=1772760 2499280 1 180 $X=1758900 $Y=2498878
X406 123 174 166 5145 4 2 5168 ADDFX2 $T=1778700 2479120 1 0 $X=1778698 $Y=2473680
X407 130 169 5145 5158 4 2 5223 ADDFX2 $T=1778700 2489200 0 0 $X=1778698 $Y=2488798
X408 5168 5155 5075 5132 4 2 5105 ADDFX2 $T=1793220 2499280 0 180 $X=1779360 $Y=2493840
X409 3606 3586 2 4 76 XNOR2X1 $T=1362240 2499280 1 180 $X=1356960 $Y=2498878
X410 3862 3865 2 4 88 XNOR2X1 $T=1428900 2499280 0 0 $X=1428898 $Y=2498878
X411 3930 3900 2 4 89 XNOR2X1 $T=1448040 2539600 0 180 $X=1442760 $Y=2534160
X412 3921 3922 2 4 3904 XNOR2X1 $T=1450680 2489200 0 180 $X=1445400 $Y=2483760
X413 3990 3989 2 4 3974 XNOR2X1 $T=1458600 2489200 0 180 $X=1453320 $Y=2483760
X414 4050 4049 2 4 97 XNOR2X1 $T=1474440 2519440 1 180 $X=1469160 $Y=2519038
X415 171 4893 2 4 4907 XNOR2X1 $T=1702140 2438800 0 0 $X=1702138 $Y=2438398
X416 4919 4920 2 4 4937 XNOR2X1 $T=1710060 2438800 0 0 $X=1710058 $Y=2438398
X417 185 5422 2 4 5443 XNOR2X1 $T=1855920 2428720 1 0 $X=1855918 $Y=2423280
X418 183 5457 2 4 5487 XNOR2X1 $T=1863840 2479120 1 0 $X=1863838 $Y=2473680
X419 5490 5486 2 4 189 XNOR2X1 $T=1874400 2418640 1 180 $X=1869120 $Y=2418238
X420 186 5488 2 4 5686 XNOR2X1 $T=1871760 2489200 0 0 $X=1871758 $Y=2488798
X421 5504 5526 2 4 5505 XNOR2X1 $T=1882980 2529520 1 180 $X=1877700 $Y=2529118
X422 5450 5561 2 4 5634 XNOR2X1 $T=1890900 2499280 0 0 $X=1890898 $Y=2498878
X423 5927 5886 2 4 203 XNOR2X1 $T=1991880 2428720 1 0 $X=1991878 $Y=2423280
X424 145 4440 127 4 2 4591 ADDHXL $T=1613040 2458960 1 0 $X=1613038 $Y=2453520
X425 126 5027 156 4 2 5062 ADDHXL $T=1760220 2479120 0 180 $X=1752960 $Y=2473680
X426 127 5087 162 4 2 5155 ADDHXL $T=1761540 2489200 1 0 $X=1761538 $Y=2483760
X427 128 5315 174 4 2 5366 ADDHXL $T=1829520 2479120 0 0 $X=1829518 $Y=2478718
X428 153 151 155 2 4 4703 XOR3X2 $T=1640100 2418640 0 0 $X=1640098 $Y=2418238
X429 5411 5335 4 5336 2 5306 AOI21XL $T=1832820 2519440 1 180 $X=1830180 $Y=2519038
X430 5331 5511 4 5540 2 5541 AOI21XL $T=1884960 2509360 0 0 $X=1884958 $Y=2508958
X431 5260 5533 4 5564 2 5585 AOI21XL $T=1892880 2448880 0 0 $X=1892878 $Y=2448478
X432 4018 3676 4046 2 4049 4 OAI2BB1X1 $T=1471140 2529520 1 0 $X=1471138 $Y=2524080
X433 4067 3996 4051 2 4080 4 OAI2BB1X1 $T=1477740 2549680 0 0 $X=1477738 $Y=2549278
X434 4093 3676 4105 2 4223 4 OAI2BB1X1 $T=1486980 2529520 0 0 $X=1486978 $Y=2529118
X435 4661 4658 4678 2 150 4 OAI2BB1X1 $T=1650000 2559760 0 180 $X=1646700 $Y=2554320
X436 5567 5549 5563 2 5560 4 OAI2BB1X1 $T=1894860 2529520 0 180 $X=1891560 $Y=2524080
X437 5804 200 5807 2 5886 4 OAI2BB1X1 $T=1954260 2428720 1 0 $X=1954258 $Y=2423280
X438 5871 5808 5841 2 5829 4 OAI2BB1X1 $T=1972740 2458960 1 180 $X=1969440 $Y=2458558
X439 3530 2 3540 4 3515 NAND2BXL $T=1349040 2428720 1 180 $X=1346400 $Y=2428318
X440 3604 2 3593 4 3505 NAND2BXL $T=1359600 2438800 0 180 $X=1356960 $Y=2433360
X441 3789 2 3770 4 3768 NAND2BXL $T=1402500 2469040 0 180 $X=1399860 $Y=2463600
X442 4106 2 4109 4 4087 NAND2BXL $T=1490280 2479120 1 180 $X=1487640 $Y=2478718
X443 4111 2 4170 4 4171 NAND2BXL $T=1503480 2479120 1 0 $X=1503478 $Y=2473680
X444 4249 2 4220 4 4134 NAND2BXL $T=1519980 2438800 0 180 $X=1517340 $Y=2433360
X445 4188 2 4203 4 4256 NAND2BXL $T=1534500 2549680 1 180 $X=1531860 $Y=2549278
X446 167 2 168 4 4919 NAND2BXL $T=1710060 2428720 1 0 $X=1710058 $Y=2423280
X447 5090 2 5088 4 5086 NAND2BXL $T=1764840 2519440 0 180 $X=1762200 $Y=2514000
X448 5117 2 5116 4 5144 NAND2BXL $T=1783320 2519440 0 0 $X=1783318 $Y=2519038
X449 5253 2 5281 4 5504 NAND2BXL $T=1861200 2529520 0 0 $X=1861198 $Y=2529118
X450 5697 2 5733 4 5718 NAND2BXL $T=1939740 2479120 1 180 $X=1937100 $Y=2478718
X451 5831 2 5841 4 5870 NAND2BXL $T=1979340 2458960 1 180 $X=1976700 $Y=2458558
X452 5900 2 5899 4 5927 NAND2BXL $T=1992540 2428720 0 0 $X=1992538 $Y=2428318
X453 128 124 4383 4343 4 2 4312 ADDFHX1 $T=1578060 2418640 1 180 $X=1562880 $Y=2418238
X454 123 126 130 4441 4 2 4402 ADDFHX1 $T=1566840 2428720 0 0 $X=1566838 $Y=2428318
X455 132 4401 4402 4395 4 2 4319 ADDFHX1 $T=1582020 2448880 0 180 $X=1566840 $Y=2443440
X456 4468 139 4454 2 138 4 AOI2BB1X2 $T=1600500 2569840 1 180 $X=1595880 $Y=2569438
X457 4404 4 4295 2 CLKINVX3 $T=1568820 2509360 0 0 $X=1568818 $Y=2508958
X458 6504 4 6460 2 CLKINVX3 $T=2152260 2428720 0 0 $X=2152258 $Y=2428318
X459 99 97 98 4 2 OR2X4 $T=1469820 2418640 0 180 $X=1465860 $Y=2413200
X460 3654 79 3662 2 4 3676 OAI2BB1X4 $T=1376760 2418640 0 0 $X=1376758 $Y=2418238
X461 2781 54 2 4 INVX8 $T=1197900 2418640 0 0 $X=1197898 $Y=2418238
X462 3676 3585 2 4 INVX8 $T=1382040 2469040 0 180 $X=1378080 $Y=2463600
X463 117 114 4239 4266 4 2 OAI2BB1X2 $T=1537140 2418640 1 180 $X=1532520 $Y=2418238
X464 210 6377 6378 6504 4 2 OAI2BB1X2 $T=2114640 2428720 0 0 $X=2114638 $Y=2428318
X465 155 151 157 4 159 2 160 4743 AOI221X1 $T=1654620 2418640 1 0 $X=1654618 $Y=2413200
X466 3716 3875 2 4 3841 3839 AOI2BB1X1 $T=1427580 2539600 0 180 $X=1424280 $Y=2534160
X467 5637 5821 2 4 5808 5805 AOI2BB1X1 $T=1957560 2458960 1 180 $X=1954260 $Y=2458558
X468 4556 4269 136 4 2 4577 OR3XL $T=1609740 2569840 0 0 $X=1609738 $Y=2569438
X469 167 170 116 2 4855 4 4893 OAI31X1 $T=1701480 2428720 1 180 $X=1697520 $Y=2428318
X470 159 2 164 4 4757 4761 NAND3XL $T=1666500 2418640 1 0 $X=1666498 $Y=2413200
X471 4048 2 116 4 CLKINVX8 $T=1536480 2448880 0 180 $X=1532520 $Y=2443440
X472 4032 3986 4 2 4081 NOR2BX4 $T=1471800 2489200 1 0 $X=1471798 $Y=2483760
X473 5303 5281 5302 2 5300 4 5296 5297 5262 OAI222XL $T=1824240 2509360 0 180 $X=1818960 $Y=2503920
X474 4202 4 2 4290 BUFX8 $T=1510740 2509360 1 0 $X=1510738 $Y=2503920
X475 4290 4 2 193 BUFX8 $T=1901460 2438800 0 0 $X=1901458 $Y=2438398
X476 4810 4773 168 4761 2 4 4855 AND4X2 $T=1684320 2428720 1 0 $X=1684318 $Y=2423280
.ENDS
***************************************
.SUBCKT ICV_55 1 3 62 64 65 67 69 70 71 73 75 77 78 80 81 83 84 1316 1317
** N=31461 EP=19 IP=95 FDC=0
X0 5439 3 5399 1 65 NAND2X1 $T=1578720 2579920 0 180 $X=1576740 $Y=2574480
X1 70 3 5439 1 5379 NAND2X1 $T=1589280 2590000 0 180 $X=1587300 $Y=2584560
X2 5399 3 73 1 5530 NAND2X1 $T=1610400 2579920 1 0 $X=1610398 $Y=2574480
X3 75 3 5585 1 5623 NAND2X1 $T=1617660 2579920 0 0 $X=1617658 $Y=2579518
X4 83 3 84 1 70 NAND2X1 $T=1651980 2590000 1 0 $X=1651978 $Y=2584560
X5 67 3 1 5439 INVX1 $T=1591260 2579920 1 180 $X=1589940 $Y=2579518
X6 69 3 1 5399 INVX1 $T=1595220 2579920 1 0 $X=1595218 $Y=2574480
X7 70 3 1 71 INVX1 $T=1597860 2579920 0 0 $X=1597858 $Y=2579518
X8 5530 3 1 5585 INVX1 $T=1605780 2579920 0 0 $X=1605778 $Y=2579518
X9 84 83 3 1 67 NOR2X2 $T=1651980 2579920 0 0 $X=1651978 $Y=2579518
X10 5623 5645 5644 3 1 NAND2X2 $T=1632840 2579920 1 180 $X=1629540 $Y=2579518
X11 78 73 1 80 5645 3 AOI21X1 $T=1634160 2579920 1 0 $X=1634158 $Y=2574480
X12 81 5644 77 3 1 XNOR2X4 $T=1636800 2590000 1 180 $X=1625580 $Y=2589598
X13 5379 64 1 3 62 XNOR2X2 $T=1576080 2590000 0 180 $X=1568820 $Y=2584560
.ENDS
***************************************
.SUBCKT ICV_54
** N=20878 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_53
** N=26494 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_52 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
** N=65 EP=40 IP=100 FDC=0
X0 3 22 PDIDGZ $T=743425 3289640 0 180 $X=715745 $Y=3104640
X1 4 23 PDIDGZ $T=823200 3289640 0 180 $X=795520 $Y=3104640
X2 5 24 PDIDGZ $T=902975 3289640 0 180 $X=875295 $Y=3104640
X3 6 25 PDIDGZ $T=982750 3289640 0 180 $X=955070 $Y=3104640
X4 7 26 PDIDGZ $T=1142300 3289640 0 180 $X=1114620 $Y=3104640
X5 8 27 PDIDGZ $T=1222075 3289640 0 180 $X=1194395 $Y=3104640
X6 9 28 PDIDGZ $T=1301845 3289640 0 180 $X=1274165 $Y=3104640
X7 10 29 PDIDGZ $T=1381615 3289640 0 180 $X=1353935 $Y=3104640
X8 11 30 PDIDGZ $T=1461385 3289640 0 180 $X=1433705 $Y=3104640
X9 12 31 PDIDGZ $T=1541155 3289640 0 180 $X=1513475 $Y=3104640
X10 13 32 PDIDGZ $T=1620925 3289640 0 180 $X=1593245 $Y=3104640
X11 14 33 PDIDGZ $T=1780465 3289640 0 180 $X=1752785 $Y=3104640
X12 15 34 PDIDGZ $T=1940005 3289640 0 180 $X=1912325 $Y=3104640
X13 16 35 PDIDGZ $T=2019775 3289640 0 180 $X=1992095 $Y=3104640
X14 17 36 PDIDGZ $T=2099545 3289640 0 180 $X=2071865 $Y=3104640
X15 18 37 PDIDGZ $T=2179320 3289640 0 180 $X=2151640 $Y=3104640
X16 19 38 PDIDGZ $T=2259095 3289640 0 180 $X=2231415 $Y=3104640
X17 20 39 PDIDGZ $T=2338870 3289640 0 180 $X=2311190 $Y=3104640
X18 21 40 PDIDGZ $T=2498420 3289640 0 180 $X=2470740 $Y=3104640
.ENDS
***************************************
.SUBCKT ICV_51 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=15 FDC=0
X3 1 5 PDO12CDG $T=2627970 0 0 0 $X=2630288 $Y=598
X4 2 4 PDO12CDG $T=2707745 0 0 0 $X=2710063 $Y=598
X5 3 6 PDO12CDG $T=2787520 0 0 0 $X=2789838 $Y=598
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=15 FDC=0
X0 1 4 PDIDGZ $T=2657970 3289640 0 180 $X=2630290 $Y=3104640
X1 2 5 PDIDGZ $T=2737745 3289640 0 180 $X=2710065 $Y=3104640
X2 3 6 PDIDGZ $T=2817520 3289640 0 180 $X=2789840 $Y=3104640
.ENDS
***************************************
.SUBCKT ICV_50
** N=2640 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_49
** N=2632 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_48
** N=2190 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_47
** N=2934 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_46
** N=1893 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_45 1 3 60 61 306 307
** N=3883 EP=6 IP=6 FDC=0
X0 61 60 3 1 INVX8 $T=2674980 1229200 1 180 $X=2671020 $Y=1228798
.ENDS
***************************************
.SUBCKT ICV_44
** N=2289 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_43 1 3 4 5 6 29 30 31 32 33 34 35 36 37 38 197 198
** N=2110 EP=17 IP=64 FDC=0
X0 203 1 30 29 3 31 OAI21XL $T=2632740 1773520 0 0 $X=2632738 $Y=1773118
X1 33 1 209 226 3 203 OAI21XL $T=2640660 1743280 0 0 $X=2640658 $Y=1742878
X2 4 1 3 35 INVX1 $T=2636040 1632400 0 0 $X=2636038 $Y=1631998
X3 6 1 3 5 INVX1 $T=2636040 1642480 1 0 $X=2636038 $Y=1637040
X4 32 1 3 209 INVX1 $T=2636040 1743280 1 0 $X=2636038 $Y=1737840
X5 30 37 1 3 221 OR2X2 $T=2645940 1773520 0 180 $X=2643300 $Y=1768080
X6 203 3 1 38 INVXL $T=2649240 1773520 0 0 $X=2649238 $Y=1773118
X7 209 33 36 1 226 3 OAI2BB1X1 $T=2635380 1753360 1 0 $X=2635378 $Y=1747920
X8 30 37 3 221 203 34 1 AOI22X1 $T=2640000 1773520 0 180 $X=2636700 $Y=1768080
.ENDS
***************************************
.SUBCKT ICV_42 1 3 4 5 36 37 38 39 40 183 184
** N=2628 EP=11 IP=21 FDC=0
X0 4 5 3 1 36 OR2XL $T=2630760 1793680 0 0 $X=2630758 $Y=1793278
X1 40 211 37 3 1 XNOR2X4 $T=2649240 1793680 1 180 $X=2638020 $Y=1793278
X2 39 38 1 3 211 XOR2X2 $T=2646600 1783600 1 180 $X=2640000 $Y=1783198
.ENDS
***************************************
.SUBCKT ICV_41
** N=3008 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40
** N=2213 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_39
** N=2169 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=2933 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_37
** N=1979 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36
** N=2474 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34 1 2 3 4
** N=13 EP=4 IP=7 FDC=0
X3 1 2 PDO12CDG $T=2947070 0 0 0 $X=2949388 $Y=598
.ENDS
***************************************
.SUBCKT ICV_33
** N=4301 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=4867 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=3877 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=5207 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=3543 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28
** N=6754 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27
** N=4184 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=3700 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=4704 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=5464 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=4068 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=3658 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=5291 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=3549 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=4282 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4
** N=13 EP=4 IP=7 FDC=0
X0 1 2 PDIDGZ $T=2977070 3289640 0 180 $X=2949390 $Y=3104640
.ENDS
***************************************
.SUBCKT ICV_17
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X2 2 4 PDO12CDG $T=3291620 234720 0 90 $X=3106620 $Y=237038
X3 1 3 PDO12CDG $T=3291620 314440 0 90 $X=3106620 $Y=316758
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X2 1 4 PDO12CDG $T=3291620 394160 0 90 $X=3106620 $Y=396478
X3 2 3 PDO12CDG $T=3291620 473880 0 90 $X=3106620 $Y=476198
.ENDS
***************************************
.SUBCKT ICV_14 1 3 4 5 6 7
** N=11 EP=6 IP=11 FDC=0
X3 1 4 PDO12CDG $T=3291620 553600 0 90 $X=3106620 $Y=555918
X4 3 5 PDO12CDG $T=3291620 713040 0 90 $X=3106620 $Y=715358
.ENDS
***************************************
.SUBCKT ICV_13 2 3 4 5 6 7
** N=12 EP=6 IP=11 FDC=0
X3 3 5 PDO12CDG $T=3291620 872480 0 90 $X=3106620 $Y=874798
X4 2 4 PDO12CDG $T=3291620 952200 0 90 $X=3106620 $Y=954518
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X2 1 4 PDO12CDG $T=3291620 1031920 0 90 $X=3106620 $Y=1034238
X3 2 3 PDO12CDG $T=3291620 1111640 0 90 $X=3106620 $Y=1113958
.ENDS
***************************************
.SUBCKT ICV_11 2 4 5 6
** N=15 EP=4 IP=7 FDC=0
X3 2 4 PDO12CDG $T=3291620 1271080 0 90 $X=3106620 $Y=1273398
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=15 FDC=0
X3 1 4 PDO12CDG $T=3291620 1430520 0 90 $X=3106620 $Y=1432838
X4 2 6 PDO12CDG $T=3291620 1510240 0 90 $X=3106620 $Y=1512558
X5 3 5 PDO12CDG $T=3291620 1589960 0 90 $X=3106620 $Y=1592278
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X2 2 4 PDO12CDG $T=3291620 1669680 0 90 $X=3106620 $Y=1671998
X3 1 3 PDO12CDG $T=3291620 1749400 0 90 $X=3106620 $Y=1751718
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=0
X2 1 4 PDO12CDG $T=3291620 1829120 0 90 $X=3106620 $Y=1831438
X3 2 3 PDO12CDG $T=3291620 1908840 0 90 $X=3106620 $Y=1911158
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4 5 6
** N=10 EP=6 IP=11 FDC=0
X3 1 3 PDO12CDG $T=3291620 1988560 0 90 $X=3106620 $Y=1990878
X4 2 4 PDO12CDG $T=3291620 2148000 0 90 $X=3106620 $Y=2150318
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=15 FDC=0
X3 1 4 PDO12CDG $T=3291620 2227720 0 90 $X=3106620 $Y=2230038
X4 2 6 PDO12CDG $T=3291620 2307440 0 90 $X=3106620 $Y=2309758
X5 3 5 PDO12CDG $T=3291620 2387160 0 90 $X=3106620 $Y=2389478
.ENDS
***************************************
.SUBCKT ICV_5 2 3 4 5
** N=9 EP=4 IP=6 FDC=0
X2 2 3 PDO12CDG $T=3291620 2546600 0 90 $X=3106620 $Y=2548918
.ENDS
***************************************
.SUBCKT ICV_4 2 3 4 5 6 7
** N=12 EP=6 IP=11 FDC=0
X3 3 4 PDO12CDG $T=3291620 2706040 0 90 $X=3106620 $Y=2708358
X4 2 5 PDO12CDG $T=3291620 2785760 0 90 $X=3106620 $Y=2788078
.ENDS
***************************************
.SUBCKT ICV_3
** N=6 EP=0 IP=1 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4
** N=9 EP=4 IP=6 FDC=0
X2 1 2 PDO12CDG $T=3291620 2945200 0 90 $X=3106620 $Y=2947518
.ENDS
***************************************
.SUBCKT ICV_1
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CHIP VDD VSS cdata_rd[4] cdata_rd[5] cdata_rd[6] cdata_rd[7] cdata_rd[8] cdata_rd[9] cdata_rd[10] cdata_rd[11] cdata_rd[12] cdata_rd[13] cdata_rd[14] cdata_rd[15] cdata_rd[16] cdata_rd[17] cdata_rd[18] cdata_rd[19] SCAN_IN SCAN_EN
+ SCAN_OUT busy iaddr[0] iaddr[1] iaddr[2] iaddr[3] iaddr[4] iaddr[5] iaddr[6] iaddr[7] iaddr[8] clk reset iaddr[9] iaddr[10] iaddr[11] ready idata[0] cwr caddr_wr[0]
+ caddr_wr[1] caddr_wr[2] caddr_wr[3] caddr_wr[4] caddr_wr[5] caddr_wr[6] caddr_wr[7] caddr_wr[8] caddr_wr[9] caddr_wr[10] caddr_wr[11] cdata_wr[0] cdata_wr[1] cdata_wr[2] cdata_wr[3] cdata_wr[4] idata[1] idata[2] idata[3] idata[4]
+ idata[5] idata[6] idata[7] idata[8] idata[9] idata[10] idata[11] idata[12] idata[13] idata[14] idata[15] idata[16] idata[17] idata[18] idata[19] cdata_wr[5] cdata_wr[6] cdata_wr[7] cdata_rd[0] cdata_rd[1]
+ cdata_rd[2] cdata_wr[8] cdata_rd[3] cdata_wr[9] cdata_wr[10] cdata_wr[11] cdata_wr[12] cdata_wr[13] cdata_wr[14] cdata_wr[15] cdata_wr[16] cdata_wr[17] cdata_wr[18] cdata_wr[19] crd caddr_rd[0] caddr_rd[1] caddr_rd[2] caddr_rd[3] caddr_rd[4]
+ caddr_rd[5] caddr_rd[6] caddr_rd[7] caddr_rd[8] caddr_rd[9] caddr_rd[10] caddr_rd[11] csel[0] csel[1] csel[2]
** N=17065 EP=110 IP=35832 FDC=0
X1 1 2 cdata_rd[4] cdata_rd[5] 17064 17065 ICV_118 $T=0 0 0 0 $X=598 $Y=185000
X2 3 4 cdata_rd[6] cdata_rd[7] 17064 17065 ICV_117 $T=0 0 0 0 $X=598 $Y=342100
X3 5 6 cdata_rd[8] cdata_rd[9] 17064 17065 ICV_116 $T=0 0 0 0 $X=598 $Y=540100
X4 8 10 cdata_rd[10] cdata_rd[11] 17064 17065 ICV_115 $T=0 0 0 0 $X=598 $Y=740700
X5 10927 10928 cdata_rd[12] cdata_rd[13] 17064 17065 ICV_114 $T=0 0 0 0 $X=598 $Y=979900
X6 11 12 cdata_rd[14] cdata_rd[15] 17064 17065 ICV_113 $T=0 0 0 0 $X=598 $Y=1139300
X7 13 14 10929 cdata_rd[16] cdata_rd[17] cdata_rd[18] 17064 17065 ICV_112 $T=0 0 0 0 $X=598 $Y=1417020
X8 15 cdata_rd[19] 17064 17065 ICV_111 $T=0 0 0 0 $X=598 $Y=1617700
X9 16 SCAN_IN 17064 17065 ICV_110 $T=0 0 0 0 $X=598 $Y=1777100
X10 10930 3479 SCAN_EN SCAN_OUT 17064 17065 ICV_109 $T=0 0 0 0 $X=598 $Y=1975060
X11 4961 253 busy iaddr[0] 17064 17065 ICV_108 $T=0 0 0 0 $X=598 $Y=2214220
X12 17 4927 iaddr[1] iaddr[2] 17064 17065 ICV_107 $T=0 0 0 0 $X=598 $Y=2414900
X13 18 19 5779 iaddr[3] iaddr[5] iaddr[4] 17064 17065 ICV_106 $T=0 0 0 0 $X=598 $Y=2574300
X15 20 iaddr[6] 17064 17065 ICV_104 $T=0 0 0 0 $X=598 $Y=2931700
X17 2247 2248 iaddr[8] iaddr[7] 17064 17065 ICV_102 $T=0 0 0 0 $X=185000 $Y=598
X30 VSS VDD 2442 2349 2366 17064 17065 ICV_89 $T=0 0 0 0 $X=185000 $Y=2574300
X33 11603 2442 clk reset 17064 17065 ICV_86 $T=0 0 0 0 $X=185000 $Y=3104600
X34 2492 4651 3479 iaddr[10] iaddr[11] iaddr[9] 17064 17065 ICV_85 $T=0 0 0 0 $X=342200 $Y=598
X40 VDD VSS 11982 2844 2846 531 2849 2835 539 11954 2851 11961 2852 11968 476 2850 538 2854 2847 11973
+ 2859 2860 11963 526 11962 515 2857 11938 523 11979 11991 11957 2865 518 535 536 537 17064 17065
+ ICV_79 $T=0 0 0 0 $X=342200 $Y=1139300
X41 VDD VSS 2928 12029 2916 2847 12027 2835 2849 2850 2851 2857 12012 2852 2913 12024 2927 2853 2854 4433
+ 12035 2935 2938 655 2859 12010 12014 542 12036 12030 2939 12032 563 3331 623 2937 2936 12011 616 513
+ 553 12013 564 2934 544 12015 12023 554 2922 595 545 12025 552 476 567 17064 17065
+ ICV_78 $T=0 0 0 0 $X=342200 $Y=1430398
X42 VSS VDD 3007 2835 3001 3008 3004 3005 2913 3006 3009 2846 2936 3020 2844 3011 2916 568 3027 3021
+ 3023 2928 2927 570 3024 2934 607 563 2935 615 655 2938 12098 12097 12088 12094 623 616 2939 577
+ 595 590 17064 17065
+ ICV_77 $T=0 0 0 0 $X=342200 $Y=1616880
X43 VDD VSS 3001 2912 3006 3005 3008 3009 3004 3011 576 568 2922 3020 3023 599 619 620 2938 3061
+ 2937 615 3021 12158 607 12155 3027 655 623 2935 12156 3068 12132 598 12157 614 612 601 563 12145
+ 617 2939 616 12144 592 12139 595 622 5657 618 621 17064 17065
+ ICV_76 $T=0 0 0 0 $X=342200 $Y=1777100
X44 VSS VDD 3061 655 615 17064 17065 ICV_75 $T=0 0 0 0 $X=342200 $Y=1990900
X50 3042 3097 ready idata[0] 17064 17065 ICV_69 $T=0 0 0 0 $X=342200 $Y=3104600
X51 VSS VDD 523 526 535 536 515 537 11963 11957 538 539 2865 11962 11973 3331 2849 11954 11991 2853
+ 518 11968 3336 3351 531 3370 3343 3341 3360 11982 3334 11961 513 3353 3354 3415 3368 3376 3411 1423
+ 3388 3371 3393 3383 3384 3385 3405 3387 3395 3397 3410 3400 3403 3399 3401 3406 3418 3413 3408 3422
+ 3407 3421 3419 3424 3427 3426 11938 11979 3453 3457 3456 3460 3458 3459 3469 3472 3478 3481 3483 3724
+ 3484 3512 3482 3487 3486 3531 3540 3488 3500 3721 3490 3504 3494 3497 3496 3542 3506 3516 3508 3511
+ 3539 3513 3514 3510 3509 3521 3522 3523 3524 3528 3525 3526 3527 3529 3530 3517 3534 3533 3536 3537
+ 3541 3548 1424 3557 3559 3560 3561 3562 3586 3563 3566 3569 3565 3571 3570 3579 3596 3714 3572 3580
+ 3601 3573 1429 3613 3578 3577 3581 3576 3584 3623 3652 3593 3587 4607 3594 3634 3574 3602 3589 3622
+ 3600 3690 3599 3669 3603 3614 3605 3665 1427 3635 3606 3610 3624 3626 3687 3618 3619 3621 3620 3650
+ 3625 3673 3632 3636 3638 3629 3640 3639 3641 3642 3644 3645 3647 1426 798 3646 1425 3653 3661 3651
+ 3649 3659 3658 3660 3668 3667 3663 3666 3670 3672 3615 3681 3675 3676 3677 3679 3609 3750 3685 3754
+ 3686 3747 3688 1428 3689 3694 3696 3740 3695 3706 3701 3756 3703 3711 3762 3717 1311 3715 3752 3730
+ 3719 3709 3760 3726 3797 3728 3738 3698 3648 3575 3725 3744 3748 3805 3755 3766 3758 3759 3763 3765
+ 3768 3775 3777 3776 3778 3779 3784 3782 3783 3781 3787 3789 3788 3792 3791 3793 3802 3790 3798 3799
+ 3796 3800 3815 3806 3808 3813 3823 1430 3827 3833 3834 15342 3835 3836 3930 15343 1431 3841 4053 3843
+ 3844 15328 3856 3846 3847 3853 3858 3863 3865 3842 3884 3878 3873 3876 3879 12464 3889 3886 3888 3895
+ 3892 3908 3890 3891 3898 3909 3900 3901 3899 3902 3903 3905 3906 3910 3912 3911 3920 3915 3916 3871
+ 3919 3918 4009 3979 3954 3950 3922 3923 3977 3985 3924 3925 3948 3693 4041 4035 3995 3928 5106 3929
+ 4010 3984 3971 3942 3970 4022 3981 3983 4016 3936 3938 4024 3969 3939 3926 3934 3947 5980 3949 3956
+ 3935 1432 3951 3952 4052 3987 3955 3957 15349 3964 4058 3960 3962 3958 3966 3967 3959 3968 4046 3972
+ 3973 3974 3975 15350 3965 6011 3982 1433 3986 3988 3999 4057 15357 15364 3993 15363 3992 3996 3998 3997
+ 823 1407 4000 15351 4002 4003 1395 4014 4012 4015 4017 4018 4020 4021 4026 4013 4027 4030 4028 4031
+ 4032 4036 4045 1258 4039 4042 4043 4056 4048 4049 4051 1245 1434 4054 4055 1281 4060 4061 4062 4068
+ 4069 4064 4065 4075 5182 4067 5134 4050 4047 4070 4236 4063 4079 4227 4078 4071 4092 4093 4223 4091
+ 4097 4098 4096 4088 4100 4120 4082 4111 4110 4090 4168 4108 4104 4107 4112 4109 4130 4118 4117 1435
+ 4174 4144 4129 4124 4133 4159 4184 4143 4128 4136 4205 4125 4137 4127 4170 4196 4132 4131 4134 4138
+ 4234 4126 4142 4139 4145 4140 1436 4151 4152 4150 4155 4153 4158 4166 4172 4169 4162 4163 4171 4167
+ 1437 4173 4175 4176 4177 4180 4179 4182 4183 4187 4188 4034 4206 4194 4198 4199 1342 4228 4210 4212
+ 4225 4230 4237 1438 4238 4242 4246 4243 4244 4245 4265 4256 4257 4259 4261 4260 4269 4270 4262 4272
+ 4282 4281 1439 4289 4300 4302 4303 4304 4305 4307 4308 4310 4320 4321 4328 1440 1441 4323 4357 4334
+ 4332 4331 4333 4335 12471 4337 4339 4346 4350 4342 1442 4351 4349 4353 4359 4365 4367 4369 4373 4370
+ 4376 4394 4372 4375 4379 4377 4378 4381 4382 4383 4384 4385 4386 4388 4390 4387 4393 4397 4399 4402
+ 4293 1443 4404 4405 17064 17065
+ ICV_62 $T=0 0 0 0 $X=660660 $Y=1138078
X52 VDD 570 VSS 4433 12088 590 12098 577 2938 2937 595 4448 623 563 4439 12097 4558 4449 4459 4461
+ 4462 4464 4471 4467 4469 4476 4501 4473 4474 4475 4477 4479 4481 4559 4485 4489 4490 4491 4496 4500
+ 4503 4504 4527 4520 4539 4525 4534 4518 12519 4530 4531 4519 861 3407 4529 3418 4532 4533 3711 3403
+ 3717 3694 4545 3413 4540 4542 4541 3419 4528 12094 4483 4551 4605 4560 4561 4566 4587 615 4569 4572
+ 4574 4579 4580 2492 3479 3589 2247 2248 3594 4607 616 4603 4933 4970 4606 253 2939 4609 4613 4943
+ 4615 4621 4626 4577 4632 4619 4591 4635 3530 3529 4651 3526 869 4641 4653 4646 4647 4655 4652 4669
+ 3548 4658 4660 4920 4817 4663 3651 4664 4662 4657 3533 4673 4676 4671 4543 4667 4677 873 4683 3578
+ 1429 4690 4687 4686 4689 3623 3580 3570 4694 3576 4696 3587 3679 4704 4714 4729 4706 3621 4708 4707
+ 4709 4710 4711 5886 4787 4715 3599 4747 3609 3615 4728 15377 10 4731 4733 4734 4735 4611 4745 4
+ 10928 15 4742 4743 4744 4746 4754 3614 6 4770 4749 4748 5 4750 8 3645 4752 3571 5084 4832
+ 3635 5049 3 4741 3622 4769 4756 5037 4759 3642 4763 4757 5061 5222 4762 4869 4941 4765 4764 4766
+ 4768 3638 4701 4794 4777 4873 3681 4778 4779 2935 3572 4782 4784 4795 4813 4781 4722 4783 2 3677
+ 4790 4785 4789 4786 3673 4828 3652 4800 1 4796 3661 4630 4797 4798 4802 4820 4805 4808 4811 4818
+ 5029 4823 3690 4814 5009 4815 4824 10788 4822 4825 10013 4717 4758 4936 4833 4834 5034 4788 4835 3714
+ 4852 4840 4849 4850 4847 4853 4855 4826 4866 4871 15378 4872 5022 4878 4879 4884 4885 4868 15350 4614
+ 4899 4897 4898 3763 4914 4902 4851 4912 4946 4907 4910 3775 4612 4917 4911 4921 4923 4926 4927 4961
+ 4950 4924 4929 4931 4934 4939 4959 4945 4957 2349 4951 2366 4952 4954 4982 4955 4956 4991 4962 4964
+ 4965 4968 4966 4969 4971 4974 4983 4976 4979 4987 4981 4984 5021 4985 5045 4993 5023 4990 4992 4997
+ 5000 4995 4998 4999 5001 5003 5004 5007 5008 5018 5012 5013 12555 5030 5042 5016 5017 3861 5019 3859
+ 5024 5028 5031 5032 5070 5040 5039 5041 903 5051 5052 5054 5056 5062 5058 5065 5090 5071 3726 5072
+ 5085 5086 5087 5088 5089 5096 3975 975 12612 5102 3967 5103 4096 5113 5180 1789 5135 3950 5120 5131
+ 5156 5117 3971 5133 5123 5125 5127 3977 4109 5128 5130 5139 5215 5136 5134 15387 5132 5144 5138 3954
+ 5140 5178 5142 4091 4118 5141 5146 3928 5150 3985 5151 5153 3992 5137 4051 5152 12586 5228 5155 5189
+ 5157 5169 5159 5161 5160 5162 4063 5188 4097 907 5173 5393 15389 5388 3942 15388 4887 4908 3984 5397
+ 4918 4050 5391 5403 5167 5408 5171 4856 5170 5193 5165 5168 12587 5172 5174 4055 4067 5191 5389 5182
+ 5366 5175 5185 5202 5181 5190 5195 5197 5198 4144 5203 5201 5200 4034 5204 909 5192 4159 5209 4378
+ 4827 5298 5216 5235 5234 5233 5454 5307 5217 5521 5230 5196 5237 5238 4760 5240 5242 5245 5248 5253
+ 5325 5251 5499 5252 5254 5255 5256 5573 5475 5359 5266 5273 5275 5278 5289 5291 5296 5304 5305 5313
+ 5306 5310 5309 4142 5315 5321 5316 5334 5328 5336 5330 5332 5347 5338 5345 5343 5344 5348 5350 5353
+ 5357 5369 5381 5382 5439 5387 5394 5429 5413 5400 5402 5406 5407 5410 5425 5421 5428 5367 5432 5447
+ 5437 5450 5441 5478 5448 5445 5451 5455 5459 5444 5462 12589 5530 5467 5464 5470 5473 5471 5472 5469
+ 5488 5477 5480 942 5491 5492 5494 5500 5501 5505 5489 5504 5507 5510 5515 5513 5512 5514 5516 5542
+ 5535 5560 5538 5540 5541 5543 4394 5545 5554 5561 5558 5564 5562 5563 5566 5575 5570 5572 5574 5576
+ 5577 5584 5585 5596 5597 5598 5602 5615 5605 5594 949 5607 12631 5617 5616 5622 5623 1990 5627 5628
+ 5629 971 5631 5632 12638 5612 5635 5638 952 983 10223 5630 979 951 966 982 953 17064 17065
+ ICV_60 $T=0 0 0 0 $X=660660 $Y=1616880
X53 VDD VSS 612 614 615 616 617 623 12156 2938 595 601 4448 598 599 12145 592 607 2939 3024
+ 12139 2937 4483 12157 4439 5670 12155 12144 5671 12158 4558 5657 5702 12132 4449 5701 5664 5665 4461 4459
+ 5666 5724 4476 3007 5676 4474 4473 4481 5677 5683 4503 4485 5697 4489 5694 5688 5687 5691 4500 4491
+ 4496 5692 4490 5690 4504 4501 5695 4520 4525 4531 5703 4527 5704 5705 861 4534 4541 4540 3711 4543
+ 3717 4528 4551 4533 4532 4561 4574 4577 4587 4591 4609 4607 5717 16 2366 20 3594 3589 253 4635
+ 17 4606 5779 5056 4614 4612 19 4619 4621 18 5024 5054 4722 4630 4811 869 4641 5785 4646 4624
+ 4647 5070 4652 4653 4654 4655 4662 5771 5751 4656 4658 4664 4602 3651 5754 4701 4661 4671 5755 3724
+ 873 4672 4617 4668 4669 4836 5791 4634 4774 4677 4683 4684 4690 5759 4778 4687 4673 3525 5764 5767
+ 4637 4694 5766 4696 3533 5772 4704 5768 3528 4707 4710 4579 4786 5784 4715 4695 4706 4714 4729 4739
+ 5800 5787 4676 4744 4815 5789 4908 4918 5788 3694 5790 5847 4758 4748 4797 5792 3658 5801 5795 4775
+ 5802 4784 8077 4780 4781 4776 5803 4788 5804 4792 5805 5814 3580 4801 5809 5810 3721 5812 5811 4806
+ 5815 15378 11603 5813 4814 5819 5822 5826 4826 4825 3488 4842 5825 5824 4835 5833 4840 5831 5877 5834
+ 4847 4887 4848 5871 4851 5913 4849 5837 5838 4855 4856 4860 5839 5964 4862 4864 4866 4868 4871 5850
+ 5844 5845 5846 4879 4880 4881 4603 5851 5852 4888 4924 5857 5855 4965 4902 5870 5867 4907 5863 5864
+ 4911 4912 4914 5866 5875 4927 5848 4921 4920 4926 4923 4928 5873 4933 4929 4931 5872 4946 5884 4934
+ 5032 5878 13659 5879 5874 5880 4937 5891 4939 5882 5888 4943 4949 4945 5883 5887 3042 4917 4948 5885
+ 4951 5890 4950 5898 4952 5892 4953 4960 4823 4959 4968 5897 4983 4966 15382 5899 4969 5905 4970 4971
+ 5896 5900 4974 3813 5910 5908 3815 5914 5924 4984 5909 5911 5912 4990 5008 4993 4992 4964 5904 5915
+ 5916 3823 3827 5001 5919 3833 4981 3837 3836 5086 5019 15343 15342 5933 5022 5021 4998 5931 5034 5029
+ 5009 5039 5936 4798 5040 903 5113 5049 5051 6067 5096 5937 5198 5942 5058 5062 5065 5949 5943 5945
+ 5195 5072 15350 5071 5947 5087 5935 5952 1656 5088 12712 4956 1559 5097 5121 5951 5958 4010 5960 5959
+ 5957 5961 5102 3979 3915 5948 5967 3954 3925 5968 3950 5120 5969 5965 5963 5950 3928 5160 5128 3948
+ 5971 3934 5973 5979 5091 5978 5974 3924 6081 5975 3971 15388 5129 15387 5132 5136 5117 6092 5131 6065
+ 4096 5169 5133 15389 5134 5178 5886 5137 6097 5138 5143 5141 5142 5981 4750 5145 5983 5146 5972 5984
+ 3955 5147 5149 6082 5986 6032 4769 5152 5153 5990 4742 5987 5991 4091 5154 3973 907 5157 3938 6050
+ 5993 3976 4802 5161 5162 5164 6047 5998 5165 6000 5061 4097 4795 5171 5174 5175 3968 4941 6005 5140
+ 4016 3936 5197 5185 6010 5941 5181 6045 5200 6012 6068 6018 4785 5201 5203 6031 5190 5191 5192 6022
+ 5204 4144 5389 909 5216 6025 4066 6027 5310 5234 6029 5230 6034 6035 6036 6037 5240 6039 6054 5256
+ 6046 5238 6048 6049 6051 5275 5297 6058 5278 6057 5289 6059 6061 5296 15412 5298 6066 6069 6063 5305
+ 5304 6072 6071 6070 5307 5253 6078 6080 5315 5316 6084 5319 6085 6086 5325 5328 5332 6091 6093 6095
+ 6098 6075 5353 5173 5359 5366 5369 5391 6118 6113 5193 6103 6114 5408 5155 6116 5381 6117 5441 5388
+ 5397 6120 5393 6125 5403 5406 6128 5455 5425 5430 5429 6134 6135 6019 6136 5413 6138 5447 5450 6139
+ 6140 6144 6145 6123 6146 5467 12711 5470 5472 5480 6151 6152 5494 942 6154 6155 5488 6156 6157 5492
+ 5500 6024 5504 5507 6167 5510 6168 5515 5516 5513 5512 6173 6174 5540 5535 5541 5538 6184 6185 6186
+ 5543 4321 4323 6188 5545 5554 6189 5563 4335 6196 5562 6194 6195 6198 6197 5574 4351 5577 4343 6203
+ 5585 4357 6207 5570 6208 5598 6209 6211 5602 5597 949 4366 6218 4359 6227 6226 6225 4381 6232 6235
+ 6228 5615 5616 6229 5622 5623 4375 5631 4379 5628 5629 6233 6234 6238 984 978 983 981 982 17064
+ 17065
+ ICV_59 $T=0 0 0 0 $X=660660 $Y=1777100
X54 15328 6239 15418 15420 6240 15423 6241 6453 6242 15428 6243 15431 15433 15357 3999 15363 15364 6244 cwr caddr_wr[1]
+ caddr_wr[3] caddr_wr[4] caddr_wr[8] caddr_wr[10] caddr_wr[11] cdata_wr[0] cdata_wr[2] cdata_wr[4] caddr_wr[0] caddr_wr[2] caddr_wr[5] caddr_wr[6] caddr_wr[7] caddr_wr[9] cdata_wr[1] cdata_wr[3] 17064 17065
+ ICV_68 $T=0 0 0 0 $X=661300 $Y=598
X57 VDD VSS 7198 7200 7201 7197 7199 7221 7222 3760 7223 7224 7227 7235 7237 7238 7243 7247 7250 7251
+ 7249 7256 7259 7283 7275 7288 7277 7274 7272 7280 7273 7276 7279 7284 7285 7286 7287 7339 17064 17065
+ ICV_65 $T=0 0 0 0 $X=661300 $Y=555900
X58 VDD VSS 1293 7526 7529 7528 7530 7527 7531 3566 7537 7538 7541 3478 3481 7542 3593 3569 7555 3575
+ 7569 7567 3618 3592 7574 3584 3625 7571 3596 3600 3645 7583 3574 3579 7585 7586 7588 3577 7587 7589
+ 3613 7590 3720 7595 7604 7602 7603 7606 7608 7609 7612 7613 7596 7631 7627 7198 7200 7197 7199 7201
+ 7645 3410 3716 3715 3718 7221 7259 7223 3709 7224 3738 3752 3754 7650 7651 3725 3762 1311 3756 3740
+ 3760 3750 3747 3728 1312 7652 7653 7222 7654 7655 7227 7658 7237 7235 7238 7250 7251 7247 7243 7249
+ 7665 1314 7666 1315 7667 7668 7256 1316 1317 7669 7286 6241 7273 7274 15420 7272 15418 3853 7275 7276
+ 7277 6240 3916 3844 4053 7279 7280 1320 7673 7670 15423 6239 7671 3876 7672 7283 7284 7674 7676 7285
+ 7675 6453 3886 7681 7288 15344 7680 1321 7679 7682 6242 7683 3905 3909 1324 7685 7686 15428 6243 15433
+ 15431 7700 7701 7705 4002 4000 7713 7715 7714 4017 7716 7720 7728 7724 7725 7339 4048 7287 4093 4068
+ 4071 4075 4082 4088 4090 7738 7740 1329 7752 7741 7763 4236 7758 4227 7754 4199 7756 7757 1338 7773
+ 7760 4184 7759 7761 7769 7772 1342 7771 7770 1340 7774 4168 7775 7779 7778 7780 7782 7783 7784 7781
+ 1339 1325 1306 1318 1330 1341 1313 1319 1323 1322 17064 17065
+ ICV_64 $T=0 0 0 0 $X=661300 $Y=739920
X59 VDD VSS 3368 3371 3369 3370 3385 3383 3384 3336 3415 3426 3424 3427 1293 7526 7527 7529 3453 7528
+ 7530 7531 3593 3458 3456 3460 7537 7538 3482 3487 7541 3484 7542 3523 3486 3497 3494 3496 3500 7555
+ 3506 3513 3516 3511 3521 3527 3536 3541 7567 7569 3563 7571 3566 3629 3613 7574 3618 3584 3581 3592
+ 3586 3600 3562 3574 3569 3645 3565 3614 3622 3571 3572 3575 3577 3623 7588 3579 7585 7583 7586 3595
+ 3601 7587 7589 7590 3596 3650 7602 3620 3610 7595 7596 3649 7603 7604 7608 7606 3652 3634 7609 3636
+ 3641 7613 7612 1306 3661 3644 3659 3647 3670 3667 3668 798 7627 7631 3685 3686 3688 3695 7651 3706
+ 3716 3715 7645 1311 3698 3752 3738 3730 3717 3709 3728 3750 3747 7650 7654 3740 3748 7652 3725 7653
+ 3756 3754 3758 3760 3762 7655 7658 1313 3759 3781 7665 3782 3777 3798 1314 7666 3797 3800 7667 7668
+ 3806 3808 3835 3834 3837 7669 3841 3847 3846 7670 3861 1319 3862 3857 1320 7671 3860 7673 7676 7672
+ 3876 3842 3853 7674 7675 3844 4053 3878 3859 7679 3888 3892 7680 3889 7681 7686 3896 1323 1324 7683
+ 1322 7682 3901 3899 3905 3909 7685 3912 3920 3930 3918 3919 3923 3922 3949 7701 1325 3956 3959 7700
+ 3962 3965 3970 7713 3976 3981 3975 3983 6487 6486 6244 4052 4057 4058 3986 3988 4046 4045 3990 3967
+ 3996 4005 7705 4009 10012 7714 4013 4015 4017 7716 7715 4020 4022 4021 4025 7720 4032 4035 4038 7724
+ 1258 4039 1024 4041 1234 4043 4042 10459 3995 4054 7728 5221 10478 7725 4066 4061 4062 4065 1245 4079
+ 4081 7738 1329 4104 4107 4110 7740 1330 4112 7741 4117 4168 4120 7774 4133 4125 4126 4128 4131 4137
+ 4139 4140 4155 4143 4145 4150 4174 7754 7752 4151 4162 4163 4223 1338 4169 7756 7757 4171 4173 7759
+ 7760 7761 4175 7763 4177 4176 7769 4184 7770 4170 7771 4236 7772 4199 7773 7775 4196 4227 1341 4206
+ 7778 7784 7780 4205 7779 7781 7758 1342 7783 7782 4234 4228 4230 4244 4245 4260 4262 4269 4272 4281
+ 4293 4393 4384 4300 4302 4369 4349 4333 4337 4343 4342 4366 4370 4372 4376 4386 4377 17064 17065
+ ICV_63 $T=0 0 0 0 $X=661300 $Y=979900
X60 VSS VDD 542 544 564 12025 12013 552 12010 545 12024 2939 563 2865 12027 567 2938 12036 2860 616
+ 623 2935 554 553 2916 12035 12032 655 12023 607 3334 12014 12029 576 3459 12011 12030 3341 4467 2912
+ 3343 12012 4462 4464 4469 12015 3351 4471 3353 3354 4477 3360 4611 3369 3376 4479 3384 1423 3387 3388
+ 3701 4545 3395 3403 3393 4540 4518 3400 3401 4519 3397 3399 4532 3408 3406 4529 3410 3694 4530 3405
+ 4528 3413 3419 3407 3640 3421 4533 3418 3422 4539 4542 4475 4560 4559 4566 4569 3457 4572 595 3472
+ 3469 4734 3589 3483 4580 3490 4602 4605 3594 4607 3411 4617 4615 3504 3508 4656 4624 3510 4613 4604
+ 3509 4654 3512 3514 4672 4626 3517 3605 3524 3488 3537 4632 3522 4665 4634 4637 3529 3525 3534 3528
+ 3531 3533 3539 4685 3540 4651 3542 4708 4662 4684 4657 4660 4661 4663 4842 4668 4667 3560 1424 3559
+ 3557 3561 4676 3572 3632 3639 3573 4686 1429 4689 3576 4695 3646 3718 1425 3602 4749 3665 4704 3669
+ 4706 3603 4709 3579 3577 4714 1427 4711 4834 4717 4856 15377 4918 3596 4747 3600 3569 3716 3606 4847
+ 3626 3613 3615 4728 14 4733 4887 3636 4735 3619 3624 4789 4683 3853 11 4741 4746 4739 4745 10927
+ 3844 4754 5061 3689 3595 4756 4752 4760 4759 5196 3629 4764 3601 3618 4908 4757 4768 4763 4731 4762
+ 4766 1426 3648 4669 3651 3653 4813 4774 12 4770 3681 3649 4779 4776 4777 4783 3666 4780 4782 3660
+ 3663 4652 3677 1428 3675 4775 4673 10929 4787 3625 3676 4792 3672 3623 3693 3580 4800 4806 4808 5183
+ 3687 4832 4801 13 5199 4817 3593 3592 4820 4825 4823 4828 4796 4851 3696 4822 4743 3698 4827 3719
+ 3720 3709 3584 4722 3703 12555 4838 5211 4836 15350 4848 4794 4872 4880 3725 4850 3575 3728 4860 4862
+ 4878 4853 4881 3755 4884 4885 3766 4888 4898 3765 4897 4899 3790 3776 3778 3863 4910 3783 4928 3784
+ 3779 4937 3787 4936 3788 3793 3789 15382 4948 3792 3796 4949 4864 3791 4954 4953 4957 3799 4961 3879
+ 3884 3802 3768 3805 4985 4960 4976 4979 4955 4982 4987 5013 4997 5023 5004 5018 3859 4999 5000 4866
+ 5003 3856 1430 5007 3860 4917 3862 4962 4991 5012 3861 5130 5016 4995 3865 1431 5091 5017 3842 5028
+ 3843 15344 5030 11603 5031 4053 3857 5041 5045 5042 3858 3896 5052 3873 3910 3871 3900 3878 3876 3895
+ 3890 3898 3891 5086 5089 5090 3744 3908 3902 3903 1445 3906 1461 5097 4612 5032 13299 5103 1803 13987
+ 3967 3975 1789 3919 4096 3929 3935 5127 5121 5123 3925 5128 3942 3951 5155 4012 3950 3952 3948 1432
+ 5135 3964 5140 3954 5151 5139 3939 5145 5143 3957 3958 5134 5147 3928 5149 4109 3971 5156 5188 3972
+ 5170 4118 5154 4051 3982 5129 3969 5144 3977 4063 3979 5167 3984 1433 4097 5168 3985 4055 3987 5164
+ 3938 5393 5172 3990 4014 5175 3997 4050 3993 5161 5182 3924 5189 5180 4016 5202 4010 5120 5200 4018
+ 3936 5201 4025 5096 4028 5193 4034 4024 4027 4060 5190 4030 4031 4124 4067 5150 5235 4127 5204 4049
+ 4047 1434 5576 4144 5197 5217 4056 4159 5215 5233 4138 5584 5228 5237 5232 4070 5223 5382 5236 4078
+ 5242 4081 5245 4064 5561 5252 5243 5255 5254 4092 5564 4098 5209 4394 5266 4100 5269 5270 5273 4108
+ 5280 4111 1435 4130 4129 5241 5297 5291 4136 4134 4132 5306 5309 1436 5313 5319 5321 4153 4152 5357
+ 4158 5334 5336 5338 4166 5341 4167 5347 5344 5343 5348 1437 4172 5350 5351 5354 4179 4180 4183 4182
+ 5367 4187 4188 4194 4198 5394 5384 5413 5387 5402 5400 4212 4210 5407 5410 5411 5421 4243 4225 5427
+ 5430 5428 1438 5439 5448 5437 5438 4237 5445 5444 5451 4242 5454 5332 5459 5462 5471 5464 4256 4257
+ 4259 4261 5469 5473 5477 5475 5478 5325 4265 4308 5489 5491 5499 5501 5505 1439 4289 5521 4303 5359
+ 5514 4304 4307 4310 5530 4378 5542 4320 4328 5572 1440 5558 4331 4332 5560 4334 4390 5566 4339 1441
+ 5607 5573 5575 4346 1442 4350 4353 5596 5594 4365 4367 4373 5605 5612 5632 4382 4387 4383 4385 4388
+ 5617 4397 4399 5627 5630 4402 4405 4404 1443 5635 5643 5638 10223 17064 17065
+ ICV_61 $T=0 0 0 0 $X=661300 $Y=1430398
X61 VSS VDD 7895 623 5666 5665 5664 5701 615 4439 5670 595 2937 4448 5671 607 7897 7896 4483 5676
+ 5677 2938 7898 655 2939 7899 2935 616 13304 5683 4558 4604 7901 7900 5692 5687 7902 5688 7904 7903
+ 5690 5697 5691 7908 5702 5705 5694 5695 7922 5724 5768 5703 5704 7923 7924 10930 5717 7925 7932 7931
+ 7933 7930 7935 7936 7937 7942 7943 7945 4611 1496 7955 5751 3651 7960 7962 5754 7964 4673 4669 4658
+ 4668 7956 3529 5785 5755 3528 4774 5771 3724 7963 7968 4664 7973 7961 7975 5759 3533 5772 5791 4701
+ 7972 7971 7976 7977 5766 7979 4695 7978 7974 5764 4848 5831 4836 5822 7981 5767 7984 4685 7986 7996
+ 7993 7992 8001 7995 4607 4860 4842 4665 5784 8006 8007 4684 5779 8008 8009 5788 5787 5790 4742 5878
+ 5789 4731 8011 8010 4750 4748 5792 4769 8033 8019 8018 8020 4941 8022 1510 8023 8105 4795 5886 8110
+ 5800 5061 4785 8034 5801 8028 8029 8181 8031 5803 5864 8035 8089 4765 8036 5805 5804 5809 15378 4802
+ 5810 4790 15519 8086 8040 5811 5812 5814 5802 5815 5870 5826 8046 5819 5825 8047 4818 5029 8048 4805
+ 5813 8114 5958 8051 8050 4824 5824 8076 4798 8057 8059 5834 8060 5833 8066 8109 5838 5837 5839 8091
+ 3097 4852 8070 4833 8084 8074 5846 5844 8077 5851 8075 4873 5847 8090 5848 5845 5795 5850 8079 8083
+ 5898 5852 4781 8082 5855 5857 5863 5892 5871 5913 5879 8268 5866 5919 5867 8096 5872 5873 5880 5874
+ 5875 5877 4869 8100 5931 8099 5882 8129 5883 5884 5885 5888 8107 5887 8115 5890 5891 5899 5897 5908
+ 5896 5113 8185 5900 8116 5904 8151 8117 8120 5909 8128 5905 8127 5910 8108 5911 8126 5912 5914 5915
+ 5916 8134 8139 8132 5085 8131 8146 8175 8148 8135 5961 4998 15523 8133 5933 8183 8165 8147 8145 4823
+ 5037 8616 8154 5935 8176 5937 8159 5960 5941 5942 5943 5121 5951 8166 5945 5049 5965 8138 5947 5948
+ 5950 5952 6012 5084 8172 8182 5973 8178 5998 5957 5968 5959 3911 4760 5963 4856 5964 5967 5106 4918
+ 5969 5924 4847 8186 4887 3926 8190 8188 8202 4851 8199 8187 4908 8189 4838 5971 5972 8222 8184 5974
+ 5125 5975 15528 6010 8233 5978 5159 8225 8231 8197 5980 8235 5981 5984 5199 8214 5983 6000 3947 8339
+ 4827 5987 15349 3960 8203 5196 5990 5211 5222 5183 5993 3974 5991 8207 8208 5986 3966 8211 8212 8217
+ 6005 6011 10013 10788 8095 4003 8226 8228 8227 8229 4026 6168 8232 4021 4036 4038 8236 8106 8237 8238
+ 4005 8245 6018 6019 15351 8247 6024 5269 8246 8224 6022 6025 8218 5221 6173 8220 5223 8253 8257 6027
+ 5243 5432 8250 6032 6031 6029 8260 5236 8243 8261 6034 5241 6035 6136 6036 6037 8263 5248 1526 8265
+ 5251 8264 8266 6039 8267 5270 15412 6048 6046 8270 6047 6050 6068 6045 6051 8274 6049 6057 6069 6054
+ 6058 6059 8280 6061 6063 6082 6065 6066 6075 8285 6072 6070 6071 8289 6078 6080 8294 6086 8293 6084
+ 5146 6085 6081 1534 8295 6095 8296 6092 6093 6091 6097 6098 8299 5341 8303 5351 8300 5354 6103 8302
+ 6128 5366 8304 6113 5389 8311 5388 6116 6117 6120 5384 6114 6118 6123 6125 8323 5411 6152 5427 5188
+ 5430 8334 6134 5438 6135 6138 4238 5189 8337 6139 6140 6144 6145 6146 6157 8346 4246 8352 6154 6151
+ 4270 8356 6155 6156 8357 8358 8361 4282 6167 6174 8366 8367 8368 4305 8374 6184 6185 6186 8375 6188
+ 8382 6189 8383 8384 6194 8386 8389 6195 8387 6196 6198 6197 1551 8390 6203 8393 8392 6207 1552 6209
+ 6211 8395 6218 8400 6228 6227 6225 6226 8403 6229 8407 6232 8405 6234 6235 6233 6238 1535 1484 1493
+ 1533 1485 1511 1483 1497 1547 1509 1481 1482 17064 17065
+ ICV_58 $T=0 0 0 0 $X=661300 $Y=1989840
X62 VDD VSS 7895 1481 7899 595 7896 7897 1482 7898 655 2938 2935 616 623 4604 2939 1483 1484 7901
+ 7902 7903 7904 1485 7908 7900 7924 7922 7923 607 1493 7925 7935 7931 7932 7936 7937 7942 7933 1496
+ 7943 4611 1497 7945 7930 7960 7956 7955 8564 7962 8475 7961 8476 7963 7964 7968 7976 7971 7972 7973
+ 8471 7974 8472 7975 8474 8473 7979 7984 7978 7981 7977 7986 7995 7992 7993 8482 7996 8007 8001 8009
+ 8490 8492 8006 8491 8008 8010 8493 8496 8011 8020 8018 8019 8022 8023 8029 8028 8031 8511 8033 8034
+ 8512 8513 8036 8514 8516 8040 8515 8521 8523 8228 4842 8524 8046 8525 8526 5822 8529 8503 8532 8060
+ 8057 8533 8212 8534 8066 8211 8535 8536 8537 8236 8217 8077 8074 8539 8109 8076 8089 8541 8232 8079
+ 8082 1509 8543 8083 8096 8086 8546 1510 8091 8084 8146 8114 8549 8550 8551 8553 8090 5864 8107 8555
+ 8127 8557 8558 8095 8559 8560 5878 8552 5848 8562 8563 8099 8571 8105 8106 8108 8182 5879 8110 8573
+ 8572 8586 1511 8172 8116 8583 8584 8576 8585 8117 8120 8587 8129 8131 8595 8132 8115 8134 8596 8133
+ 8135 8138 8139 8175 8154 8601 8145 8147 5931 8605 8606 8148 8604 8151 8652 8622 8181 8159 8613 8614
+ 8615 5847 8619 8621 8165 8618 8623 8633 5891 8635 8629 8628 8616 8186 5871 5877 8634 8128 8188 8184
+ 8183 5913 8639 8203 8640 8185 5964 8126 8187 8645 8190 8689 5987 6000 5979 8197 8199 5972 8189 8202
+ 8659 8662 5983 8663 8176 8207 8208 8665 5991 8668 8669 8656 8218 8673 8220 5978 8675 8224 8671 8226
+ 8227 8229 8681 8686 8237 8238 8698 8693 8699 8688 8243 8245 8246 8247 8694 8250 8257 5232 8253 8166
+ 8263 8260 8708 8261 1526 8264 8710 8265 8266 8267 8268 8270 5280 8274 8771 8280 8723 8730 8285 8289
+ 1533 8293 8728 1535 8729 8294 8296 8295 8731 5330 8732 8733 8299 5345 8738 8300 8742 8743 8303 8304
+ 8744 8745 8748 8746 8747 8311 8323 8334 8214 8337 8346 8352 8356 8357 8358 8361 8789 1547 8367 8366
+ 8368 8374 8375 8382 8383 8384 8395 8386 8387 8389 1551 8390 8392 1552 6208 8393 8400 8403 8405 8407
+ 17064 17065
+ ICV_57 $T=0 0 0 0 $X=661300 $Y=2230000
X63 VSS VDD 8471 8473 8472 8474 8475 8476 8482 8490 8492 8493 8496 8491 8503 8511 8512 8513 8514 8515
+ 8516 8521 8523 8524 8525 8526 8051 8059 8532 8533 8529 8535 8534 8537 8536 8543 8539 8541 8546 8550
+ 8549 8551 8552 8553 8555 8990 8557 8558 8559 8560 8563 8562 8564 8572 8571 8573 8576 8583 8585 8584
+ 8586 8606 8604 8587 8595 9004 8120 8596 8134 8138 8616 8993 8175 8129 8176 8994 8996 8601 8997 8995
+ 8184 8605 8133 9000 8154 5978 8139 9005 9006 9007 8614 8629 8613 9009 8615 8187 8618 8115 8621 8619
+ 9011 8197 9013 8622 9017 8202 8635 8628 6000 8633 8634 8135 8639 8214 8640 8645 8652 8623 8656 8659
+ 8663 8665 8203 8668 8208 8207 8669 8671 8673 8675 8681 8723 8698 8688 8689 8693 8694 8686 8699 8708
+ 8662 8710 8728 8729 8733 8730 8731 8732 8738 8742 8743 8302 8747 8745 8746 8744 8748 8771 8789 17064
+ 17065
+ ICV_56 $T=0 0 0 0 $X=661300 $Y=2413200
X64 VDD VSS 8990 8994 8993 8995 8996 9011 8997 9006 9000 9004 9005 9007 9017 9009 9013 17064 17065 ICV_55 $T=0 0 0 0 $X=661300 $Y=2574300
X67 8047 8070 8050 8048 15519 8035 8075 5113 8100 5085 15523 8178 8225 8233 8222 8231 8235 8339 15528 idata[1]
+ idata[2] idata[3] idata[4] idata[5] idata[6] idata[7] idata[8] idata[9] idata[10] idata[11] idata[12] idata[13] idata[14] idata[15] idata[16] idata[17] idata[18] idata[19] 17064 17065
+ ICV_52 $T=0 0 0 0 $X=661300 $Y=3104600
X68 6487 6486 10012 cdata_wr[6] cdata_wr[5] cdata_wr[7] 17064 17065 ICV_51 $T=0 0 0 0 $X=2614470 $Y=598
X69 5034 5009 10013 cdata_rd[0] cdata_rd[1] cdata_rd[2] 17064 17065 ICV_35 $T=0 0 0 0 $X=2614470 $Y=3104600
X75 VDD VSS 12464 12471 17064 17065 ICV_45 $T=0 0 0 0 $X=2630300 $Y=1139300
X77 VSS VDD 951 952 953 978 966 1990 10223 971 12638 5643 12631 983 10262 17064 17065 ICV_43 $T=0 0 0 0 $X=2630300 $Y=1617700
X78 VDD VSS 982 983 984 12711 981 10262 966 17064 17065 ICV_42 $T=0 0 0 0 $X=2630300 $Y=1777100
X85 10459 cdata_wr[8] 17064 17065 ICV_34 $T=0 0 0 0 $X=2815200 $Y=598
X101 10788 cdata_rd[3] 17064 17065 ICV_18 $T=0 0 0 0 $X=2815200 $Y=3104600
X103 1024 10478 cdata_wr[10] cdata_wr[9] 17064 17065 ICV_16 $T=0 0 0 0 $X=3106600 $Y=185000
X104 1234 1245 cdata_wr[12] cdata_wr[11] 17064 17065 ICV_15 $T=0 0 0 0 $X=3106600 $Y=342100
X105 1258 1281 cdata_wr[13] cdata_wr[14] 17064 17065 ICV_14 $T=0 0 0 0 $X=3106600 $Y=540100
X106 1395 4069 cdata_wr[16] cdata_wr[15] 17064 17065 ICV_13 $T=0 0 0 0 $X=3106600 $Y=740700
X107 1407 3998 cdata_wr[18] cdata_wr[17] 17064 17065 ICV_12 $T=0 0 0 0 $X=3106600 $Y=979900
X108 823 cdata_wr[19] 17064 17065 ICV_11 $T=0 0 0 0 $X=3106600 $Y=1139300
X109 1445 1461 13299 crd caddr_rd[1] caddr_rd[0] 17064 17065 ICV_10 $T=0 0 0 0 $X=3106600 $Y=1417020
X110 975 12612 caddr_rd[3] caddr_rd[2] 17064 17065 ICV_9 $T=0 0 0 0 $X=3106600 $Y=1617700
X111 5102 12712 caddr_rd[5] caddr_rd[4] 17064 17065 ICV_8 $T=0 0 0 0 $X=3106600 $Y=1777100
X112 1559 5949 caddr_rd[6] caddr_rd[7] 17064 17065 ICV_7 $T=0 0 0 0 $X=3106600 $Y=1975060
X113 1656 5936 6067 caddr_rd[8] caddr_rd[10] caddr_rd[9] 17064 17065 ICV_6 $T=0 0 0 0 $X=3106600 $Y=2214220
X114 13659 caddr_rd[11] 17064 17065 ICV_5 $T=0 0 0 0 $X=3106600 $Y=2414900
X115 1803 1789 csel[0] csel[1] 17064 17065 ICV_4 $T=0 0 0 0 $X=3106600 $Y=2574300
X117 13987 csel[2] 17064 17065 ICV_2 $T=0 0 0 0 $X=3106600 $Y=2931700
.ENDS
***************************************
