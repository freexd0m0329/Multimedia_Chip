D:/Documents/Git/Multimedia_Chip/opt/Design_kit/CBDK_TSMC018_Arm_v3.2/CIC/SOCE/lef/tpb973gv_6lm.lef