// Verilog HDL NetList 
//   timeStamp 2009 10 20 13 39 9 
//   author "Avanti Corporation."
//   program "A2Hdl" 
//   design library: io_tpz973gv
//   cell name     : io_tpz973gv.CEL (version 1)
module PAD50ARU ();
endmodule
module PAD60NU ();
endmodule
module PAD70NU ();
endmodule
module PAD80NU ();
endmodule
module PDD04DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD02SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD02DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB04SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB04DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB02SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDB02DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PCORNER ();
endmodule 
module PCI66SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PCI66DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PCI33SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PCI33DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDT08DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT04DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT02DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDO24CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO16CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO12CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO08CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO04CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDO02CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PDISDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDIDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDDWDGZ ( C , PAD , REN );
    output C ;
    input PAD ;
    input REN ;
endmodule 
module PDDW24DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW16DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW12DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW08DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW04DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDW02DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDDSDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDDDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDD24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDD04SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDXOE2DG ( E , XC , XIN , XOUT );
    input E ;
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXOE1DG ( E , XC , XIN , XOUT );
    input E ;
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXO03DG ( XC , XIN , XOUT );
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXO02DG ( XC , XIN , XOUT );
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDXO01DG ( XC , XIN , XOUT );
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PDUWDGZ ( C , PAD , REN );
    output C ;
    input PAD ;
    input REN ;
endmodule 
module PDUW24DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW16DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW12DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW08DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW04DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUW02DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PDUSDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDUDGZ ( C , PAD );
    output C ;
    input PAD ;
endmodule 
module PDU24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU04SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU04DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU02SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDU02DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PDT24DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT16DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PDT12DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRO08CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PRDW24DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRDW16DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRDW12DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRDW08DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRD24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRD08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRCUT ();
endmodule 
module PRB24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRB08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PFILLER5 ();
endmodule 
module PFILLER20 ();
endmodule 
module PFILLER1 ();
endmodule 
module PFILLER10 ();
endmodule 
module PFILLER05 ();
endmodule 
module PFILLER0005 ();
endmodule 
module PDXOE3DG ( E , XC , XIN , XOUT );
    input E ;
    output XC ;
    input XIN ;
    output XOUT ;
endmodule 
module PVSS3DGZ ();
endmodule 
module PVSS2DGZ ( VSSPST );
    inout VSSPST ;
endmodule 
module PVSS2ANA ( AVSS );
    inout AVSS ;
endmodule 
module PVSS1DGZ ();
endmodule 
module PVSS1ANA ( AVSS );
    inout AVSS ;
endmodule 
module PVDD2POC ( VD33 );
    inout VD33 ;
endmodule 
module PVDD2DGZ ( VD33 );
    inout VD33 ;
endmodule 
module PVDD2ANA ( AVDD );
    inout AVDD ;
endmodule 
module PVDD1DGZ ();
endmodule 
module PVDD1ANA ( AVDD );
    inout AVDD ;
endmodule 
module PRUW24DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRUW16DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRUW12DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRUW08DGZ ( C , I , OEN , PAD , REN );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
    input REN ;
endmodule 
module PRU24SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU24DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU16SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU16DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU12SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU12DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU08SDGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRU08DGZ ( C , I , OEN , PAD );
    output C ;
    input I ;
    input OEN ;
    inout PAD ;
endmodule 
module PRT24DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRT16DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRT12DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRT08DGZ ( I , OEN , PAD );
    input I ;
    input OEN ;
    output PAD ;
endmodule 
module PRO24CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PRO16CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 
module PRO12CDG ( I , PAD );
    input I ;
    output PAD ;
endmodule 

